//: version "1.8.7"

module CPA(A1, C0, B2, A2, B3, S3, A0, B0, C4, S1, B1, S2, A3, S0);
//: interface  /sz:(223, 91) /bd:[ Ti0>B0(136/223) Ti1>A0(118/223) Ti2>B1(103/223) Ti3>A1(83/223) Ti4>B2(66/223) Ti5>A2(48/223) Ti6>B3(29/223) Ti7>A3(11/223) Ri0>C0(34/91) Lo0<C4(39/91) Bo0<S3(39/223) Bo1<S2(76/223) Bo2<S1(127/223) Bo3<S0(175/223) ]
input A0;    //: /sn:0 {0}(1242,224)(1242,281)(1246,281)(1246,291){1}
output S1;    //: /sn:0 /dp:1 {0}(960,474)(960,508)(959,508)(959,522){1}
input C0;    //: /sn:0 {0}(1483,376)(1445,376)(1445,374)(1435,374){1}
input A3;    //: /sn:0 {0}(194,240)(194,276)(195,276)(195,286){1}
input A2;    //: /sn:0 {0}(526,227)(526,272)(527,272)(527,282){1}
input B2;    //: /sn:0 {0}(633,228)(633,275)(632,275)(632,282){1}
output C4;    //: /sn:0 {0}(75,372)(117,372)(117,373)(127,373){1}
input B1;    //: /sn:0 {0}(993,203)(993,273)(995,273)(995,283){1}
output S0;    //: /sn:0 /dp:1 {0}(1316,482)(1316,529)(1318,529)(1318,540){1}
input A1;    //: /sn:0 {0}(886,204)(886,273)(890,273)(890,283){1}
input B3;    //: /sn:0 {0}(298,244)(298,276)(300,276)(300,286){1}
output S3;    //: /sn:0 {0}(266,523)(266,487)(265,487)(265,477){1}
input B0;    //: /sn:0 {0}(1347,227)(1347,281)(1351,281)(1351,291){1}
output S2;    //: /sn:0 /dp:1 {0}(597,473)(597,511)(602,511)(602,526){1}
wire w6;    //: /sn:0 {0}(1079,366)(1168,366)(1168,378)(1178,378){1}
wire w4;    //: /sn:0 {0}(716,365)(812,365)(812,370)(822,370){1}
wire w3;    //: /sn:0 {0}(384,369)(459,369){1}
//: enddecls

  //: input g4 (A1) @(886,202) /sn:0 /R:3 /w:[ 0 ]
  //: input g8 (C0) @(1485,376) /sn:0 /R:2 /w:[ 0 ]
  FA g16 (.A(A1), .B(B1), .Cin(w6), .Cout(w4), .S(S1));   //: @(823, 284) /sz:(255, 189) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  //: input g3 (B2) @(633,226) /sn:0 /R:3 /w:[ 0 ]
  FA g17 (.A(A0), .B(B0), .Cin(C0), .Cout(w6), .S(S0));   //: @(1179, 292) /sz:(255, 189) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<1 Bo0<0 ]
  //: input g2 (A2) @(526,225) /sn:0 /R:3 /w:[ 0 ]
  //: input g1 (B3) @(298,242) /sn:0 /R:3 /w:[ 0 ]
  //: output g10 (S3) @(266,520) /sn:0 /R:3 /w:[ 0 ]
  //: input g6 (A0) @(1242,222) /sn:0 /R:3 /w:[ 0 ]
  //: input g7 (B0) @(1347,225) /sn:0 /R:3 /w:[ 0 ]
  //: output g9 (C4) @(78,372) /sn:0 /R:2 /w:[ 0 ]
  //: output g12 (S1) @(959,519) /sn:0 /R:3 /w:[ 1 ]
  FA g14 (.A(A3), .B(B3), .Cin(w3), .Cout(C4), .S(S3));   //: @(128, 287) /sz:(255, 189) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<1 ]
  //: input g5 (B1) @(993,201) /sn:0 /R:3 /w:[ 0 ]
  //: output g11 (S2) @(602,523) /sn:0 /R:3 /w:[ 1 ]
  FA g15 (.A(A2), .B(B2), .Cin(w4), .Cout(w3), .S(S2));   //: @(460, 283) /sz:(255, 189) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  //: input g0 (A3) @(194,238) /sn:0 /R:3 /w:[ 0 ]
  //: output g13 (S0) @(1318,537) /sn:0 /R:3 /w:[ 1 ]

endmodule

module FA(S, Cout, Cin, B, A);
//: interface  /sz:(255, 189) /bd:[ Ti0>B(172/255) Ti1>A(67/255) Ri0>Cin(82/189) Lo0<Cout(86/189) Bo0<S(137/255) ]
input B;    //: /sn:0 {0}(171,166)(186,166)(186,140)(219,140){1}
//: {2}(223,140)(251,140){3}
//: {4}(221,142)(221,245)(392,245){5}
input A;    //: /sn:0 {0}(157,108)(185,108)(185,135)(198,135){1}
//: {2}(202,135)(251,135){3}
//: {4}(200,137)(200,240)(392,240){5}
input Cin;    //: /sn:0 {0}(182,222)(336,222)(336,188){1}
//: {2}(338,186)(348,186)(348,205)(379,205){3}
//: {4}(336,184)(336,161)(346,161){5}
output Cout;    //: /sn:0 /dp:1 {0}(476,236)(507,236)(507,213)(518,213){1}
output S;    //: /sn:0 /dp:1 {0}(367,159)(480,159)(480,152)(490,152){1}
wire w7;    //: /sn:0 {0}(413,243)(445,243)(445,238)(455,238){1}
wire w4;    //: /sn:0 {0}(400,208)(445,208)(445,233)(455,233){1}
wire w2;    //: /sn:0 {0}(272,138)(297,138){1}
//: {2}(301,138)(336,138)(336,156)(346,156){3}
//: {4}(299,140)(299,210)(379,210){5}
//: enddecls

  //: output g4 (S) @(487,152) /sn:0 /w:[ 1 ]
  and g8 (.I0(A), .I1(B), .Z(w7));   //: @(403,243) /sn:0 /delay:" 1" /w:[ 5 5 0 ]
  //: output g3 (Cout) @(515,213) /sn:0 /w:[ 1 ]
  //: input g2 (Cin) @(180,222) /sn:0 /w:[ 0 ]
  //: input g1 (B) @(169,166) /sn:0 /w:[ 0 ]
  //: joint g10 (w2) @(299, 138) /w:[ 2 -1 1 4 ]
  xor g6 (.I0(w2), .I1(Cin), .Z(S));   //: @(357,159) /sn:0 /delay:" 2" /w:[ 3 5 0 ]
  and g7 (.I0(Cin), .I1(w2), .Z(w4));   //: @(390,208) /sn:0 /delay:" 1" /w:[ 3 5 0 ]
  //: joint g9 (Cin) @(336, 186) /w:[ 2 4 -1 1 ]
  //: joint g12 (B) @(221, 140) /w:[ 2 -1 1 4 ]
  xor g5 (.I0(A), .I1(B), .Z(w2));   //: @(262,138) /sn:0 /delay:" 2" /w:[ 3 3 0 ]
  //: joint g11 (A) @(200, 135) /w:[ 2 -1 1 4 ]
  //: input g0 (A) @(155,108) /sn:0 /w:[ 0 ]
  or g13 (.I0(w4), .I1(w7), .Z(Cout));   //: @(466,236) /sn:0 /delay:" 1" /w:[ 1 1 0 ]

endmodule

module main;    //: root_module
wire w13;    //: /sn:0 {0}(248,212)(248,248)(260,248)(260,238){1}
wire w4;    //: /sn:0 {0}(312,-61)(327,-61)(327,119){1}
wire w0;    //: /sn:0 {0}(202,65)(238,65)(238,119){1}
wire w3;    //: /sn:0 {0}(277,-42)(312,-42)(312,119){1}
wire w12;    //: /sn:0 {0}(285,212)(285,249)(301,249)(301,239){1}
wire w18;    //: /sn:0 {0}(173,153)(173,159)(208,159){1}
wire w10;    //: /sn:0 {0}(384,212)(384,250)(405,250)(405,240){1}
wire w1;    //: /sn:0 {0}(236,38)(257,38)(257,119){1}
wire w8;    //: /sn:0 {0}(202,96)(220,96)(220,119){1}
wire w14;    //: /sn:0 {0}(236,9)(275,9)(275,119){1}
wire w11;    //: /sn:0 {0}(336,212)(336,249)(353,249)(353,239){1}
wire w2;    //: /sn:0 {0}(276,-14)(292,-14)(292,119){1}
wire w5;    //: /sn:0 {0}(312,-90)(345,-90)(345,119){1}
wire w9;    //: /sn:0 {0}(432,98)(442,98)(442,154)(433,154){1}
//: enddecls

  led g4 (.I(w10));   //: @(405,233) /sn:0 /w:[ 1 ] /type:0
  //: switch g8 (w0) @(185,65) /sn:0 /w:[ 0 ] /st:0
  led g3 (.I(w11));   //: @(353,232) /sn:0 /w:[ 1 ] /type:0
  led g2 (.I(w12));   //: @(301,232) /sn:0 /w:[ 1 ] /type:0
  led g1 (.I(w13));   //: @(260,231) /sn:0 /w:[ 1 ] /type:0
  //: switch g10 (w14) @(219,9) /sn:0 /w:[ 0 ] /st:0
  //: switch g6 (w9) @(415,98) /sn:0 /w:[ 0 ] /st:0
  //: switch g7 (w8) @(185,96) /sn:0 /w:[ 0 ] /st:0
  //: switch g9 (w1) @(219,38) /sn:0 /w:[ 0 ] /st:0
  //: switch g12 (w3) @(260,-42) /sn:0 /w:[ 0 ] /st:0
  led g5 (.I(w18));   //: @(173,146) /sn:0 /w:[ 0 ] /type:0
  //: switch g11 (w2) @(259,-14) /sn:0 /w:[ 0 ] /st:0
  //: switch g14 (w5) @(295,-90) /sn:0 /w:[ 0 ] /st:0
  CPA g0 (.B0(w5), .A0(w4), .B1(w3), .A1(w2), .B2(w14), .A2(w1), .B3(w0), .A3(w8), .C0(w9), .C4(w18), .S3(w13), .S2(w12), .S1(w11), .S0(w10));   //: @(209, 120) /sz:(223, 91) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Ti3>1 Ti4>1 Ti5>1 Ti6>1 Ti7>1 Ri0>1 Lo0<1 Bo0<0 Bo1<0 Bo2<0 Bo3<0 ]
  //: switch g13 (w4) @(295,-61) /sn:0 /w:[ 0 ] /st:0

endmodule
