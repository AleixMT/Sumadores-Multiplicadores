//: version "1.8.7"

module main;    //: root_module
wire w32;    //: /sn:0 {0}(302,-62)(302,-165)(252,-165){1}
wire w37;    //: /sn:0 {0}(388,-62)(388,-137)(349,-137){1}
wire w24;    //: /sn:0 {0}(246,20)(275,20){1}
wire w23;    //: /sn:0 /dp:1 {0}(272,-62)(272,-80)(254,-80){1}
wire w36;    //: /sn:0 {0}(378,-62)(378,-108)(350,-108){1}
wire [3:0] w25;    //: /sn:0 /dp:1 {0}(342,138)(342,73){1}
wire w35;    //: /sn:0 {0}(368,-62)(368,-80)(350,-80){1}
wire [3:0] w8;    //: /sn:0 {0}(299,-27)(299,-46)(287,-46)(287,-56){1}
wire w30;    //: /sn:0 {0}(292,-62)(292,-137)(253,-137){1}
wire [3:0] w22;    //: /sn:0 {0}(364,-27)(364,-46)(383,-46)(383,-56){1}
wire w27;    //: /sn:0 /dp:1 {0}(282,-62)(282,-108)(254,-108){1}
wire w33;    //: /sn:0 {0}(398,-62)(398,-165)(348,-165){1}
wire w26;    //: /sn:0 /dp:1 {0}(430,26)(399,26){1}
//: enddecls

  //: switch g28 (w27) @(237,-108) /sn:0 /w:[ 1 ] /st:1
  //: switch g27 (w23) @(237,-80) /sn:0 /w:[ 1 ] /st:1
  //: switch g32 (w36) @(333,-108) /sn:0 /w:[ 1 ] /st:1
  CLA g19 (.B(w22), .A(w8), .C0(w24), .S(w25), .C4(w26));   //: @(276, -26) /sz:(122, 98) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Bo0<1 Ro0<1 ]
  //: switch g31 (w37) @(332,-137) /sn:0 /w:[ 1 ] /st:1
  //: switch g25 (w30) @(236,-137) /sn:0 /w:[ 1 ] /st:1
  //: switch g29 (w33) @(331,-165) /sn:0 /w:[ 1 ] /st:1
  led g21 (.I(w26));   //: @(437,26) /sn:0 /R:3 /w:[ 0 ] /type:0
  concat g24 (.I0(w23), .I1(w27), .I2(w30), .I3(w32), .Z(w8));   //: @(287,-57) /sn:0 /R:3 /w:[ 0 0 0 0 1 ] /dr:0
  //: switch g23 (w24) @(229,20) /sn:0 /w:[ 0 ] /st:1
  led g22 (.I(w25));   //: @(342,145) /sn:0 /R:2 /w:[ 0 ] /type:1
  //: switch g26 (w32) @(235,-165) /sn:0 /w:[ 1 ] /st:1
  //: switch g33 (w35) @(333,-80) /sn:0 /w:[ 1 ] /st:1
  concat g30 (.I0(w35), .I1(w36), .I2(w37), .I3(w33), .Z(w22));   //: @(383,-57) /sn:0 /R:3 /w:[ 0 0 0 0 1 ] /dr:0

endmodule

module PFA(Pi, A, Ci, Gi, S, B);
//: interface  /sz:(100, 97) /bd:[ Ti0>A(14/100) Ti1>B(50/100) Li0>Ci(46/97) Bo0<Gi(61/100) Ro0<S(32/97) Ro1<Pi(67/97) ]
input B;    //: /sn:0 {0}(184,223)(195,223){1}
//: {2}(199,223)(226,223)(226,207)(234,207){3}
//: {4}(197,225)(197,256){5}
//: {6}(199,258)(308,258){7}
//: {8}(197,260)(197,293)(309,293){9}
output Gi;    //: /sn:0 /dp:1 {0}(330,291)(354,291){1}
input A;    //: /sn:0 {0}(186,202)(214,202){1}
//: {2}(218,202)(234,202){3}
//: {4}(216,204)(216,251){5}
//: {6}(218,253)(308,253){7}
//: {8}(216,255)(216,288)(309,288){9}
output Pi;    //: /sn:0 /dp:1 {0}(329,256)(351,256){1}
input Ci;    //: /sn:0 /dp:1 {0}(305,227)(274,227)(274,241)(187,241){1}
output S;    //: /sn:0 {0}(358,225)(326,225){1}
wire w11;    //: /sn:0 {0}(255,205)(295,205)(295,222)(305,222){1}
//: enddecls

  //: output g8 (Pi) @(348,256) /sn:0 /w:[ 1 ]
  //: input g4 (A) @(184,202) /sn:0 /w:[ 0 ]
  //: joint g13 (B) @(197, 258) /w:[ 6 5 -1 8 ]
  xor g3 (.I0(A), .I1(B), .Z(w11));   //: @(245,205) /sn:0 /delay:" 2" /w:[ 3 3 0 ]
  xor g2 (.I0(w11), .I1(Ci), .Z(S));   //: @(316,225) /sn:0 /delay:" 2" /w:[ 1 0 1 ]
  or g1 (.I0(A), .I1(B), .Z(Pi));   //: @(319,256) /sn:0 /w:[ 7 7 0 ]
  //: joint g11 (B) @(197, 223) /w:[ 2 -1 1 4 ]
  //: joint g10 (A) @(216, 202) /w:[ 2 -1 1 4 ]
  //: input g6 (Ci) @(185,241) /sn:0 /w:[ 1 ]
  //: output g9 (Gi) @(351,291) /sn:0 /w:[ 1 ]
  //: output g7 (S) @(355,225) /sn:0 /w:[ 0 ]
  //: input g5 (B) @(182,223) /sn:0 /w:[ 0 ]
  and g0 (.I0(A), .I1(B), .Z(Gi));   //: @(320,291) /sn:0 /w:[ 9 9 0 ]
  //: joint g12 (A) @(216, 253) /w:[ 6 5 -1 8 ]

endmodule

module CLL(P2, C0, P1, G1, G0, P3, G3, C3, G2, C2, C1, P0, C4);
//: interface  /sz:(622, 40) /bd:[ Ti0>P3(584/622) Ti1>G3(554/622) Ti2>C3(477/622) Ti3>P2(412/622) Ti4>G2(384/622) Ti5>C2(323/622) Ti6>P1(261/622) Ti7>G1(232/622) Ti8>C1(152/622) Ti9>P0(100/622) Ti10>G0(67/622) Li0>C0(19/40) To0<C0(176/622) Ro0<C4(19/40) ]
input G2;    //: /sn:0 {0}(386,5)(342,5)(342,99)(-50,99){1}
//: {2}(-52,97)(-52,-213){3}
//: {4}(-52,101)(-52,237)(240,237){5}
input C0;    //: /sn:0 {0}(118,-214)(118,-192){1}
//: {2}(120,-190)(135,-190)(135,-199)(229,-199){3}
//: {4}(118,-188)(118,-138){5}
//: {6}(120,-136)(131,-136)(131,-119)(229,-119){7}
//: {8}(118,-134)(118,-49){9}
//: {10}(120,-47)(134,-47)(134,-40)(239,-40){11}
//: {12}(118,-45)(118,134)(183,134)(183,141)(243,141){13}
input P1;    //: /sn:0 {0}(243,151)(7,151)(7,140)(-8,140){1}
//: {2}(-10,138)(-10,2){3}
//: {4}(-8,0)(103,0)(103,10)(236,10){5}
//: {6}(-10,-2)(-10,-28){7}
//: {8}(-8,-30)(239,-30){9}
//: {10}(-10,-32)(-10,-91){11}
//: {12}(-8,-93)(3,-93)(3,-71)(229,-71){13}
//: {14}(-10,-95)(-10,-115){15}
//: {16}(-8,-117)(99,-117)(99,-109)(229,-109){17}
//: {18}(-10,-119)(-10,-214){19}
//: {20}(-10,142)(-10,175)(1,175)(1,185)(240,185){21}
output C3;    //: /sn:0 {0}(407,-3)(448,-3){1}
input G0;    //: /sn:0 {0}(75,-217)(75,-155){1}
//: {2}(77,-153)(155,-153)(155,-154)(379,-154){3}
//: {4}(75,-151)(75,-78){5}
//: {6}(77,-76)(229,-76){7}
//: {8}(75,-74)(75,3){9}
//: {10}(77,5)(236,5){11}
//: {12}(75,7)(75,180)(240,180){13}
output C4;    //: /sn:0 {0}(411,192)(459,192){1}
output C2;    //: /sn:0 {0}(402,-101)(441,-101)(441,-100)(451,-100){1}
input P3;    //: /sn:0 {0}(240,223)(-112,223)(-112,214)(-121,214){1}
//: {2}(-123,212)(-123,186){3}
//: {4}(-121,184)(-112,184)(-112,195)(240,195){5}
//: {6}(-123,182)(-123,157){7}
//: {8}(-121,155)(-106,155)(-106,161)(243,161){9}
//: {10}(-123,153)(-123,-212){11}
//: {12}(-123,216)(-123,242)(240,242){13}
input G1;    //: /sn:0 {0}(381,-96)(231,-96)(231,-90)(27,-90){1}
//: {2}(25,-92)(25,-214){3}
//: {4}(25,-88)(25,27){5}
//: {6}(27,29)(39,29)(39,50)(238,50){7}
//: {8}(25,31)(25,207)(127,207)(127,213)(240,213){9}
input G3;    //: /sn:0 /dp:1 {0}(-151,-212)(-151,266)(318,266)(318,202)(390,202){1}
output C1;    //: /sn:0 {0}(400,-156)(445,-156){1}
input P0;    //: /sn:0 /dp:11 {0}(239,-35)(144,-35)(144,-32)(58,-32){1}
//: {2}(56,-34)(56,-119){3}
//: {4}(58,-121)(69,-121)(69,-114)(229,-114){5}
//: {6}(56,-123)(56,-184){7}
//: {8}(58,-186)(140,-186)(140,-194)(229,-194){9}
//: {10}(56,-188)(56,-217){11}
//: {12}(56,-30)(56,140)(73,140)(73,146)(243,146){13}
input P2;    //: /sn:0 {0}(240,190)(-67,190)(-67,177)(-76,177){1}
//: {2}(-78,175)(-78,154)(-80,154)(-80,134){3}
//: {4}(-78,132)(17,132)(17,125)(63,125)(63,156)(243,156){5}
//: {6}(-80,130)(-80,78)(-79,78)(-79,40){7}
//: {8}(-77,38)(-48,38)(-48,55)(238,55){9}
//: {10}(-77,38)(-79,38)(-79,19){11}
//: {12}(-77,17)(-65,17)(-65,15)(236,15){13}
//: {14}(-79,15)(-79,-15){15}
//: {16}(-77,-17)(60,-17)(60,-25)(239,-25){17}
//: {18}(-79,-19)(-79,-212){19}
//: {20}(-78,179)(-78,208)(60,208)(60,218)(240,218){21}
wire w14;    //: /sn:0 {0}(257,10)(378,10)(378,-5)(386,-5){1}
wire w23;    //: /sn:0 {0}(261,187)(377,187)(377,192)(390,192){1}
wire w20;    //: /sn:0 {0}(264,151)(384,151)(384,182)(390,182){1}
wire w8;    //: /sn:0 {0}(250,-73)(371,-73)(371,-101)(381,-101){1}
wire w17;    //: /sn:0 {0}(259,53)(378,53)(378,0)(386,0){1}
wire w11;    //: /sn:0 {0}(260,-33)(379,-33)(379,-10)(386,-10){1}
wire w2;    //: /sn:0 {0}(250,-196)(335,-196)(335,-159)(379,-159){1}
wire w5;    //: /sn:0 {0}(250,-114)(372,-114)(372,-106)(381,-106){1}
wire w29;    //: /sn:0 {0}(261,240)(380,240)(380,197)(390,197){1}
wire w26;    //: /sn:0 {0}(261,218)(360,218)(360,187)(390,187){1}
//: enddecls

  //: input g4 (P2) @(-79,-214) /sn:0 /R:3 /w:[ 19 ]
  //: input g8 (C0) @(118,-216) /sn:0 /R:3 /w:[ 0 ]
  and g13 (.I0(G0), .I1(P1), .I2(P2), .Z(w14));   //: @(247,10) /sn:0 /w:[ 11 5 13 0 ]
  //: joint g37 (P0) @(56, -32) /w:[ 1 2 -1 12 ]
  //: joint g34 (P1) @(-10, -93) /w:[ 12 14 -1 11 ]
  //: input g3 (P1) @(-10,-216) /sn:0 /R:3 /w:[ 19 ]
  //: input g2 (G1) @(25,-216) /sn:0 /R:3 /w:[ 3 ]
  //: input g1 (G0) @(75,-219) /sn:0 /R:3 /w:[ 0 ]
  and g11 (.I0(G0), .I1(P1), .Z(w8));   //: @(240,-73) /sn:0 /w:[ 7 13 0 ]
  and g16 (.I0(G0), .I1(P1), .I2(P2), .I3(P3), .Z(w23));   //: @(251,187) /sn:0 /w:[ 13 21 0 5 0 ]
  //: joint g28 (P0) @(56, -186) /w:[ 8 10 -1 7 ]
  //: joint g50 (P3) @(-123, 155) /w:[ 8 10 -1 7 ]
  and g10 (.I0(C0), .I1(P0), .I2(P1), .Z(w5));   //: @(240,-114) /sn:0 /w:[ 7 5 17 0 ]
  //: joint g27 (C0) @(118, -190) /w:[ 2 1 -1 4 ]
  //: joint g32 (P1) @(-10, -117) /w:[ 16 18 -1 15 ]
  or g19 (.I0(w2), .I1(G0), .Z(C1));   //: @(390,-156) /sn:0 /w:[ 1 3 0 ]
  //: joint g38 (P1) @(-10, -30) /w:[ 8 10 -1 7 ]
  //: input g6 (P3) @(-123,-214) /sn:0 /R:3 /w:[ 11 ]
  //: joint g53 (P2) @(-78, 177) /w:[ 1 2 -1 20 ]
  //: joint g57 (P3) @(-123, 214) /w:[ 1 2 -1 12 ]
  //: input g7 (G3) @(-151,-214) /sn:0 /R:3 /w:[ 0 ]
  and g9 (.I0(C0), .I1(P0), .Z(w2));   //: @(240,-196) /sn:0 /w:[ 3 9 0 ]
  and g15 (.I0(C0), .I1(P0), .I2(P1), .I3(P2), .I4(P3), .Z(w20));   //: @(254,151) /sn:0 /w:[ 13 13 0 5 9 0 ]
  or g20 (.I0(w5), .I1(w8), .I2(G1), .Z(C2));   //: @(392,-101) /sn:0 /w:[ 1 1 0 0 ]
  //: joint g31 (P0) @(56, -121) /w:[ 4 6 -1 3 ]
  //: joint g39 (P2) @(-79, -17) /w:[ 16 18 -1 15 ]
  //: joint g48 (P1) @(-10, 140) /w:[ 1 2 -1 20 ]
  //: joint g43 (G1) @(25, 29) /w:[ 6 5 -1 8 ]
  //: output g25 (C3) @(445,-3) /sn:0 /w:[ 1 ]
  //: joint g29 (G0) @(75, -153) /w:[ 2 1 -1 4 ]
  and g17 (.I0(G1), .I1(P2), .I2(P3), .Z(w26));   //: @(251,218) /sn:0 /w:[ 9 21 0 0 ]
  //: joint g42 (P2) @(-79, 17) /w:[ 12 14 -1 11 ]
  //: input g5 (G2) @(-52,-215) /sn:0 /R:3 /w:[ 3 ]
  and g14 (.I0(G1), .I1(P2), .Z(w17));   //: @(249,53) /sn:0 /w:[ 7 9 0 ]
  //: joint g44 (P2) @(-79, 38) /w:[ 8 -1 10 7 ]
  or g21 (.I0(w11), .I1(w14), .I2(w17), .I3(G2), .Z(C3));   //: @(397,-3) /sn:0 /w:[ 1 1 1 0 0 ]
  //: joint g36 (C0) @(118, -47) /w:[ 10 9 -1 12 ]
  //: output g24 (C2) @(448,-100) /sn:0 /w:[ 1 ]
  //: joint g41 (P1) @(-10, 0) /w:[ 4 6 -1 3 ]
  //: output g23 (C1) @(442,-156) /sn:0 /w:[ 1 ]
  //: joint g40 (G0) @(75, 5) /w:[ 10 9 -1 12 ]
  //: joint g54 (P3) @(-123, 184) /w:[ 4 6 -1 3 ]
  //: input g0 (P0) @(56,-219) /sn:0 /R:3 /w:[ 11 ]
  //: joint g45 (G2) @(-52, 99) /w:[ 1 2 -1 4 ]
  or g22 (.I0(w20), .I1(w26), .I2(w23), .I3(w29), .I4(G3), .Z(C4));   //: @(401,192) /sn:0 /w:[ 1 1 1 1 1 0 ]
  //: joint g35 (G1) @(25, -90) /w:[ 1 2 -1 4 ]
  //: output g26 (C4) @(456,192) /sn:0 /w:[ 1 ]
  and g12 (.I0(C0), .I1(P0), .I2(P1), .I3(P2), .Z(w11));   //: @(250,-33) /sn:0 /w:[ 11 0 9 17 0 ]
  and g18 (.I0(G2), .I1(P3), .Z(w29));   //: @(251,240) /sn:0 /w:[ 5 13 0 ]
  //: joint g33 (G0) @(75, -76) /w:[ 6 5 -1 8 ]
  //: joint g30 (C0) @(118, -136) /w:[ 6 5 -1 8 ]
  //: joint g49 (P2) @(-80, 132) /w:[ 4 6 -1 3 ]

endmodule

module CLA(A, S, C0, C4, B);
//: interface  /sz:(122, 98) /bd:[ Ti0>B[3:0](88/122) Ti1>A[3:0](23/122) Li0>C0(46/98) Bo0<S[3:0](66/122) Ro0<C4(52/98) ]
input [3:0] B;    //: /sn:0 /dp:1 {0}(40,86)(137,86){1}
//: {2}(138,86)(301,86){3}
//: {4}(302,86)(459,86){5}
//: {6}(460,86)(621,86){7}
//: {8}(622,86)(726,86){9}
input C0;    //: /sn:0 {0}(30,251)(40,251){1}
//: {2}(44,251)(52,251)(52,215)(87,215){3}
//: {4}(42,253)(42,372)(68,372){5}
input [3:0] A;    //: /sn:0 {0}(42,61)(101,61){1}
//: {2}(102,61)(138,61)(138,61)(265,61){3}
//: {4}(266,61)(423,61){5}
//: {6}(424,61)(585,61){7}
//: {8}(586,61)(732,61){9}
output C4;    //: /sn:0 {0}(739,372)(692,372){1}
output [3:0] S;    //: /sn:0 /dp:1 {0}(760,529)(739,529){1}
wire w6;    //: /sn:0 {0}(302,170)(302,90){1}
wire w7;    //: /sn:0 {0}(266,170)(266,65){1}
wire w16;    //: /sn:0 {0}(511,244)(530,244)(530,322)(488,322)(488,351){1}
wire w15;    //: /sn:0 {0}(433,269)(433,337)(441,337)(441,351){1}
wire w19;    //: /sn:0 {0}(586,173)(586,65){1}
wire w4;    //: /sn:0 /dp:1 {0}(112,267)(112,309)(113,309)(113,351){1}
wire w0;    //: /sn:0 {0}(138,168)(138,90){1}
wire w3;    //: /sn:0 /dp:1 {0}(733,534)(381,534)(381,203)(353,203){1}
wire w34;    //: /sn:0 /dp:1 {0}(556,351)(556,220)(571,220){1}
wire w21;    //: /sn:0 {0}(595,272)(595,339)(596,339)(596,351){1}
wire w31;    //: /sn:0 /dp:1 {0}(392,351)(392,217)(409,217){1}
wire w28;    //: /sn:0 {0}(236,351)(236,217)(251,217){1}
wire w20;    //: /sn:0 {0}(673,241)(690,241)(690,321)(645,321)(645,351){1}
wire w1;    //: /sn:0 {0}(102,168)(102,65){1}
wire w8;    //: /sn:0 {0}(733,524)(541,524)(541,218)(511,218){1}
wire w18;    //: /sn:0 {0}(622,173)(622,90){1}
wire w11;    //: /sn:0 /dp:1 {0}(189,236)(202,236)(202,326)(160,326)(160,351){1}
wire w2;    //: /sn:0 {0}(733,544)(212,544)(212,201)(189,201){1}
wire w12;    //: /sn:0 {0}(460,170)(460,90){1}
wire w10;    //: /sn:0 {0}(733,514)(705,514)(705,206)(673,206){1}
wire w13;    //: /sn:0 {0}(424,170)(424,65){1}
wire w5;    //: /sn:0 {0}(353,238)(371,238)(371,326)(345,326)(345,351){1}
wire w9;    //: /sn:0 {0}(278,269)(278,335)(284,335)(284,351){1}
//: enddecls

  //: input g4 (A) @(40,61) /sn:0 /w:[ 0 ]
  tran g8(.Z(w7), .I(A[1]));   //: @(266,59) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  tran g13(.Z(w18), .I(B[3]));   //: @(622,84) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  PFA g3 (.A(w19), .B(w18), .Ci(w34), .Gi(w21), .S(w10), .Pi(w20));   //: @(572, 174) /sz:(100, 97) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Bo0<0 Ro0<1 Ro1<0 ]
  PFA g2 (.A(w13), .B(w12), .Ci(w31), .Gi(w15), .S(w8), .Pi(w16));   //: @(410, 171) /sz:(100, 97) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Bo0<0 Ro0<1 Ro1<0 ]
  PFA g1 (.A(w7), .B(w6), .Ci(w28), .Gi(w9), .S(w3), .Pi(w5));   //: @(252, 171) /sz:(100, 97) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Bo0<0 Ro0<1 Ro1<0 ]
  tran g11(.Z(w12), .I(B[2]));   //: @(460,84) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  //: joint g16 (C0) @(42, 251) /w:[ 2 -1 1 4 ]
  tran g10(.Z(w13), .I(A[2]));   //: @(424,59) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  //: output g19 (S) @(757,529) /sn:0 /w:[ 0 ]
  tran g6(.Z(w1), .I(A[0]));   //: @(102,59) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  tran g9(.Z(w6), .I(B[1]));   //: @(302,84) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  tran g7(.Z(w0), .I(B[0]));   //: @(138,84) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  //: input g15 (C0) @(28,251) /sn:0 /w:[ 0 ]
  //: output g17 (C4) @(736,372) /sn:0 /w:[ 0 ]
  //: input g5 (B) @(38,86) /sn:0 /w:[ 0 ]
  CLL g14 (.P3(w20), .G3(w21), .P2(w16), .G2(w15), .P1(w5), .G1(w9), .P0(w11), .G0(w4), .C0(C0), .C3(w34), .C2(w31), .C1(w28), .C4(C4));   //: @(69, 352) /sz:(622, 43) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Ti3>1 Ti4>1 Ti5>1 Ti6>1 Ti7>1 Li0>5 To0<0 To1<0 To2<0 Ro0<1 ]
  PFA g0 (.A(w1), .B(w0), .Ci(C0), .Gi(w4), .S(w2), .Pi(w11));   //: @(88, 169) /sz:(100, 97) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>3 Bo0<0 Ro0<1 Ro1<0 ]
  tran g12(.Z(w19), .I(A[3]));   //: @(586,59) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  concat g18 (.I0(w2), .I1(w3), .I2(w8), .I3(w10), .Z(S));   //: @(738,529) /sn:0 /w:[ 0 0 0 0 1 ] /dr:0

endmodule
