//: version "1.8.7"

module CarryLookahead_Logic(C3, P0, C4, G0, P3, G1, P1, P2, PG, C1, C2, G3, Cin, GG, G2);
//: interface  /sz:(328, 96) /bd:[ Ti0>G0(286/328) Ti1>P0(267/328) Ti2>G1(210/328) Ti3>P1(189/328) Ti4>G2(139/328) Ti5>P2(117/328) Ti6>G3(55/328) Ti7>P3(28/328) Ri0>Cin(46/96) To0<C3(86/328) To1<C2(159/328) To2<C1(228/328) Lo0<Cout(39/96) Bo0<PG(276/328) Bo1<GG(313/328) ]
input G2;    //: /sn:0 /dp:1 {0}(559,261)(542,261)(542,278)(532,278)(532,309)(218,309){1}
//: {2}(214,309)(134,309)(134,313)(49,313){3}
//: {4}(216,311)(216,429)(416,429){5}
output GG;    //: /sn:0 /dp:1 {0}(550,450)(626,450)(626,415)(636,415){1}
input P1;    //: /sn:0 /dp:1 {0}(53,230)(62,230){1}
//: {2}(66,230)(89,230)(89,213)(146,213){3}
//: {4}(150,213)(331,213)(331,157)(336,157){5}
//: {6}(148,215)(148,508)(431,508){7}
//: {8}(64,232)(64,456)(230,456){9}
output C3;    //: /sn:0 /dp:1 {0}(580,259)(592,259)(592,278)(595,278){1}
//: {2}(599,278)(618,278)(618,269)(622,269){3}
//: {4}(597,280)(597,297)(617,297){5}
output PG;    //: /sn:0 /dp:1 {0}(251,458)(306,458){1}
input G0;    //: /sn:0 {0}(72,169)(218,169){1}
//: {2}(222,169)(254,169)(254,139)(264,139)(264,129){3}
//: {4}(266,127)(270,127){5}
//: {6}(262,127)(258,127){7}
//: {8}(220,171)(220,503)(431,503){9}
output C4;    //: /sn:0 /dp:1 {0}(699,317)(734,317)(734,333)(758,333){1}
output C2;    //: /sn:0 /dp:1 {0}(417,169)(429,169)(429,178)(432,178){1}
//: {2}(436,178)(454,178)(454,177)(456,177){3}
//: {4}(434,180)(434,246)(466,246){5}
input Cin;    //: /sn:0 {0}(85,65)(97,65){1}
//: {2}(101,65)(108,65){3}
//: {4}(99,67)(99,82)(151,82){5}
input P3;    //: /sn:0 {0}(40,343)(48,343)(48,323)(141,323){1}
//: {2}(145,323)(599,323)(599,302)(617,302){3}
//: {4}(143,325)(143,333){5}
//: {6}(145,335)(325,335){7}
//: {8}(329,335)(406,335)(406,424)(416,424){9}
//: {10}(327,337)(327,448)(377,448){11}
//: {12}(381,448)(417,448){13}
//: {14}(379,450)(379,493)(431,493){15}
//: {16}(143,337)(143,466)(230,466){17}
input G1;    //: /sn:0 /dp:1 {0}(396,171)(382,171)(382,180)(372,180)(372,249)(184,249){1}
//: {2}(180,249)(51,249){3}
//: {4}(182,251)(182,453)(417,453){5}
input G3;    //: /sn:0 {0}(30,372)(447,372){1}
//: {2}(451,372)(682,372)(682,339)(670,339)(670,319)(678,319){3}
//: {4}(449,374)(449,410)(487,410)(487,443)(529,443){5}
input P0;    //: /sn:0 {0}(72,145)(88,145)(88,147)(102,147){1}
//: {2}(106,147)(135,147)(135,87)(151,87){3}
//: {4}(104,149)(104,443)(186,443)(186,449){5}
//: {6}(188,451)(230,451){7}
//: {8}(184,451)(179,451){9}
output C1;    //: /sn:0 /dp:1 {0}(291,125)(295,125)(295,112)(304,112)(304,127)(314,127){1}
//: {2}(318,127)(349,127)(349,125)(352,125){3}
//: {4}(316,129)(316,152)(336,152){5}
input P2;    //: /sn:0 /dp:1 {0}(417,458)(394,458){1}
//: {2}(390,458)(342,458)(342,281)(143,281)(143,288){3}
//: {4}(145,290)(469,290)(469,283)(479,283)(479,272)(468,272)(468,266)(456,266)(456,251)(466,251){5}
//: {6}(141,290)(101,290)(101,284)(50,284){7}
//: {8}(143,292)(143,449)(187,449)(187,459){9}
//: {10}(189,461)(230,461){11}
//: {12}(185,461)(179,461){13}
//: {14}(392,460)(392,490)(421,490)(421,498)(431,498){15}
wire w6;    //: /sn:0 {0}(437,427)(447,427)(447,448)(529,448){1}
wire w7;    //: /sn:0 {0}(438,453)(529,453){1}
wire w4;    //: /sn:0 {0}(357,155)(364,155)(364,166)(396,166){1}
wire w3;    //: /sn:0 {0}(487,249)(514,249)(514,256)(559,256){1}
wire w8;    //: /sn:0 {0}(452,500)(519,500)(519,458)(529,458){1}
wire w2;    //: /sn:0 {0}(638,300)(668,300)(668,314)(678,314){1}
wire w5;    //: /sn:0 {0}(258,124)(258,118){1}
//: {2}(260,116)(265,116)(265,122)(270,122){3}
//: {4}(258,114)(258,85)(172,85){5}
//: enddecls

  or g44 (.I0(G3), .I1(w6), .I2(w7), .I3(w8), .Z(GG));   //: @(540,450) /sn:0 /tech:unit /w:[ 5 1 1 1 0 ]
  and g8 (.I0(C1), .I1(P1), .Z(w4));   //: @(347,155) /sn:0 /tech:unit /w:[ 5 5 0 ]
  and g4 (.I0(Cin), .I1(P0), .Z(w5));   //: @(162,85) /sn:0 /tech:unit /w:[ 5 3 5 ]
  //: joint g47 (G3) @(449, 372) /w:[ 2 -1 1 4 ]
  or g16 (.I0(w3), .I1(G2), .Z(C3));   //: @(570,259) /sn:0 /tech:unit /w:[ 1 0 0 ]
  or g3 (.I0(w5), .I1(G0), .Z(C1));   //: @(281,125) /sn:0 /tech:unit /w:[ 3 5 0 ]
  //: joint g26 (C1) @(316, 127) /w:[ 2 -1 1 4 ]
  //: output g17 (C3) @(619,269) /sn:0 /w:[ 3 ]
  //: input g2 (P0) @(70,145) /sn:0 /w:[ 0 ]
  //: joint g30 (P1) @(64, 230) /w:[ 2 -1 1 8 ]
  //: output g23 (C4) @(755,333) /sn:0 /w:[ 1 ]
  //: joint g39 (P3) @(327, 335) /w:[ 8 -1 7 10 ]
  //: joint g24 (Cin) @(99, 65) /w:[ 2 -1 1 4 ]
  //: input g1 (G0) @(70,169) /sn:0 /w:[ 0 ]
  and g29 (.I0(P0), .I1(P1), .I2(P2), .I3(P3), .Z(PG));   //: @(241,458) /sn:0 /tech:unit /w:[ 7 9 11 17 0 ]
  //: input g18 (P3) @(38,343) /sn:0 /w:[ 0 ]
  or g10 (.I0(w4), .I1(G1), .Z(C2));   //: @(407,169) /sn:0 /tech:unit /w:[ 1 0 0 ]
  //: joint g25 (G0) @(264, 127) /w:[ 4 -1 6 3 ]
  //: input g6 (G1) @(49,249) /sn:0 /w:[ 3 ]
  and g35 (.I0(P3), .I1(G2), .Z(w6));   //: @(427,427) /sn:0 /w:[ 9 5 0 ]
  //: joint g9 (w5) @(258, 116) /w:[ 2 4 -1 1 ]
  //: input g7 (P1) @(51,230) /sn:0 /w:[ 0 ]
  //: joint g31 (P2) @(143, 290) /w:[ 4 3 6 8 ]
  or g22 (.I0(w2), .I1(G3), .Z(C4));   //: @(689,317) /sn:0 /tech:unit /w:[ 1 3 0 ]
  //: joint g45 (P1) @(148, 213) /w:[ 4 -1 3 6 ]
  and g41 (.I0(P3), .I1(P2), .I2(G0), .I3(P1), .Z(w8));   //: @(442,500) /sn:0 /w:[ 15 15 9 7 0 ]
  //: joint g36 (P3) @(143, 335) /w:[ 6 5 -1 16 ]
  //: joint g33 (P3) @(143, 323) /w:[ 2 -1 1 4 ]
  //: joint g42 (P3) @(379, 448) /w:[ 12 -1 11 14 ]
  //: joint g40 (G1) @(182, 249) /w:[ 1 -1 2 4 ]
  //: input g12 (P2) @(48,284) /sn:0 /w:[ 7 ]
  //: joint g46 (G0) @(220, 169) /w:[ 2 -1 1 8 ]
  //: output g34 (PG) @(303,458) /sn:0 /w:[ 1 ]
  //: joint g28 (C3) @(597, 278) /w:[ 2 -1 1 4 ]
  and g14 (.I0(C2), .I1(P2), .Z(w3));   //: @(477,249) /sn:0 /tech:unit /w:[ 5 5 0 ]
  //: output g5 (C1) @(349,125) /sn:0 /w:[ 3 ]
  //: output g11 (C2) @(453,177) /sn:0 /w:[ 3 ]
  //: joint g21 (P0) @(186, 451) /w:[ 6 5 8 -1 ]
  //: input g19 (G3) @(28,372) /sn:0 /w:[ 0 ]
  //: joint g32 (P2) @(187, 461) /w:[ 10 9 12 -1 ]
  and g20 (.I0(C3), .I1(P3), .Z(w2));   //: @(628,300) /sn:0 /tech:unit /w:[ 5 3 0 ]
  //: joint g43 (P2) @(392, 458) /w:[ 1 -1 2 14 ]
  and g38 (.I0(P3), .I1(G1), .I2(P2), .Z(w7));   //: @(428,453) /sn:0 /tech:unit /w:[ 13 5 0 0 ]
  //: joint g15 (P0) @(104, 147) /w:[ 2 -1 1 4 ]
  //: input g0 (Cin) @(83,65) /sn:0 /w:[ 0 ]
  //: output g48 (GG) @(633,415) /sn:0 /w:[ 1 ]
  //: joint g27 (C2) @(434, 178) /w:[ 2 -1 1 4 ]
  //: joint g37 (G2) @(216, 309) /w:[ 1 -1 2 4 ]
  //: input g13 (G2) @(47,313) /sn:0 /w:[ 3 ]

endmodule

module main;    //: root_module
wire w6;    //: /sn:0 {0}(346,-81)(356,-81)(356,108){1}
wire w16;    //: /sn:0 {0}(272,-59)(326,-59)(326,108){1}
wire w13;    //: /sn:0 {0}(443,216)(443,206){1}
wire w7;    //: /sn:0 {0}(270,-24)(306,-24)(306,108){1}
wire w4;    //: /sn:0 {0}(390,-174)(434,-174)(434,108){1}
wire w0;    //: /sn:0 {0}(97,164)(97,174)(112,174)(112,148)(166,148){1}
wire w10;    //: /sn:0 {0}(183,-6)(284,-6)(284,108){1}
wire w8;    //: /sn:0 {0}(183,22)(253,22)(253,108){1}
wire w17;    //: /sn:0 {0}(385,-137)(395,-137)(395,108){1}
wire w14;    //: /sn:0 {0}(480,216)(480,206){1}
wire w2;    //: /sn:0 {0}(508,70)(518,70)(518,85)(506,85)(506,155)(496,155){1}
wire w11;    //: /sn:0 {0}(346,-120)(377,-120)(377,108){1}
wire w15;    //: /sn:0 {0}(174,87)(195,87)(195,108){1}
wire w5;    //: /sn:0 {0}(434,-199)(453,-199)(453,108){1}
wire w9;    //: /sn:0 {0}(179,53)(222,53)(222,108){1}
//: enddecls

  //: switch g8 (w11) @(329,-120) /sn:0 /w:[ 0 ] /st:0
  //: switch g4 (w10) @(166,-6) /sn:0 /w:[ 0 ] /st:0
  //: switch g3 (w8) @(166,22) /sn:0 /w:[ 0 ] /st:0
  //: switch g2 (w9) @(162,53) /sn:0 /w:[ 0 ] /st:0
  //: switch g1 (w15) @(157,87) /sn:0 /w:[ 0 ] /st:0
  //: switch g10 (w4) @(373,-174) /sn:0 /w:[ 0 ] /st:0
  //: switch g6 (w16) @(255,-59) /sn:0 /w:[ 0 ] /st:0
  //: switch g9 (w17) @(368,-137) /sn:0 /w:[ 0 ] /st:0
  //: switch g7 (w6) @(329,-81) /sn:0 /w:[ 0 ] /st:0
  //: switch g12 (w2) @(491,70) /sn:0 /w:[ 0 ] /st:0
  //: switch g11 (w5) @(417,-199) /sn:0 /w:[ 0 ] /st:0
  //: switch g5 (w7) @(253,-24) /sn:0 /w:[ 0 ] /st:0
  CarryLookahead_Logic g0 (.P3(w15), .G3(w9), .P2(w10), .G2(w7), .P1(w6), .G1(w11), .P0(w4), .G0(w5), .Cin(w2), .C1(w17), .C2(w16), .C3(w8), .Cout(w0), .GG(w14), .PG(w13));   //: @(167, 109) /sz:(328, 96) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Ti3>1 Ti4>1 Ti5>1 Ti6>1 Ti7>1 Ri0>1 To0<1 To1<1 To2<1 Lo0<1 Bo0<1 Bo1<1 ]
  led g13 (.I(w0));   //: @(97,157) /sn:0 /w:[ 0 ] /type:0

endmodule
