//: version "1.8.7"

module ha(S, CO, B, A);
//: interface  /sz:(55, 65) /bd:[ Li0>B(35/65) Li1>A(20/65) Ro0<CO(41/65) Ro1<S(21/65) ]
input B;    //: /sn:0 {0}(170,290)(233,290)(233,291)(292,291){1}
//: {2}(296,291)(373,291)(373,258)(377,258){3}
//: {4}(294,289)(294,259)(302,259){5}
input A;    //: /sn:0 {0}(171,218)(275,218){1}
//: {2}(279,218)(365,218)(365,253)(377,253){3}
//: {4}(277,220)(277,254)(302,254){5}
output CO;    //: /sn:0 /dp:1 {0}(323,257)(352,257){1}
output S;    //: /sn:0 {0}(428,255)(407,255)(407,256)(398,256){1}
//: enddecls

  xor g4 (.I0(A), .I1(B), .Z(S));   //: @(388,256) /sn:0 /delay:" 2" /w:[ 3 3 1 ]
  //: output g3 (S) @(425,255) /sn:0 /w:[ 0 ]
  //: output g2 (CO) @(349,257) /sn:0 /w:[ 1 ]
  //: input g1 (B) @(168,290) /sn:0 /w:[ 0 ]
  //: joint g6 (A) @(277, 218) /w:[ 2 -1 1 4 ]
  //: joint g7 (B) @(294, 291) /w:[ 2 4 1 -1 ]
  and g5 (.I0(A), .I1(B), .Z(CO));   //: @(313,257) /sn:0 /tech:unit /w:[ 5 5 0 ]
  //: input g0 (A) @(169,218) /sn:0 /w:[ 0 ]

endmodule

module RCA_4b(Z0, Y0, X3, X2, X1, Z2, Y2, Z1, Y3, Z4, Z6, Z3, Y1, Z7, X0, Z5);
//: interface  /sz:(128, 136) /bd:[ Ti0>X0(116/128) Ti1>X1(107/128) Ti2>X2(98/128) Ti3>X3(87/128) Ti4>Y0(47/128) Ti5>Y1(34/128) Ti6>Y2(25/128) Ti7>Y3(14/128) Bo0<Z0(116/128) Bo1<Z1(104/128) Bo2<Z2(92/128) Bo3<Z3(81/128) Bo4<Z4(70/128) Bo5<Z5(60/128) Bo6<Z6(51/128) Bo7<Z7(41/128) ]
input Y3;    //: /sn:0 {0}(550,279)(540,279){1}
input X1;    //: /sn:0 {0}(330,78)(330,88){1}
input Y2;    //: /sn:0 {0}(547,245)(537,245){1}
output Z0;    //: /sn:0 /dp:1 {0}(426,177)(426,367){1}
output Z3;    //: /sn:0 /dp:1 {0}(277,347)(277,357){1}
input X2;    //: /sn:0 {0}(260,80)(260,90){1}
output Z6;    //: /sn:0 /dp:1 {0}(115,342)(115,352){1}
output Z4;    //: /sn:0 /dp:1 {0}(213,344)(213,354){1}
output Z5;    //: /sn:0 /dp:1 {0}(160,346)(160,356){1}
output Z7;    //: /sn:0 /dp:1 {0}(58,344)(58,354){1}
input X0;    //: /sn:0 {0}(415,78)(415,146)(424,146)(424,156){1}
output Z2;    //: /sn:0 /dp:1 {0}(333,346)(333,356){1}
output Z1;    //: /sn:0 /dp:1 {0}(391,339)(391,349){1}
input Y0;    //: /sn:0 {0}(544,146)(429,146)(429,156){1}
input Y1;    //: /sn:0 {0}(546,197)(536,197){1}
input X3;    //: /sn:0 {0}(210,82)(210,92){1}
//: enddecls

  //: output g8 (Z0) @(426,364) /sn:0 /R:3 /w:[ 1 ]
  //: input g4 (Y0) @(546,146) /sn:0 /R:2 /w:[ 0 ]
  and g16 (.I0(Y0), .I1(X0), .Z(Z0));   //: @(426,167) /sn:0 /R:3 /w:[ 1 1 0 ]
  //: input g3 (X3) @(210,80) /sn:0 /R:3 /w:[ 0 ]
  //: input g2 (X2) @(260,78) /sn:0 /R:3 /w:[ 0 ]
  //: input g1 (X1) @(330,76) /sn:0 /R:3 /w:[ 0 ]
  //: output g10 (Z2) @(333,353) /sn:0 /R:3 /w:[ 1 ]
  //: input g6 (Y2) @(549,245) /sn:0 /R:2 /w:[ 0 ]
  //: output g9 (Z1) @(391,346) /sn:0 /R:3 /w:[ 1 ]
  //: input g7 (Y3) @(552,279) /sn:0 /R:2 /w:[ 0 ]
  //: output g12 (Z4) @(213,351) /sn:0 /R:3 /w:[ 1 ]
  //: output g14 (Z6) @(115,349) /sn:0 /R:3 /w:[ 1 ]
  //: output g11 (Z3) @(277,354) /sn:0 /R:3 /w:[ 1 ]
  //: input g5 (Y1) @(548,197) /sn:0 /R:2 /w:[ 0 ]
  //: output g15 (Z7) @(58,351) /sn:0 /R:3 /w:[ 1 ]
  //: input g0 (X0) @(415,76) /sn:0 /R:3 /w:[ 0 ]
  //: output g13 (Z5) @(160,353) /sn:0 /R:3 /w:[ 1 ]

endmodule

module FA(Cout, S, Cin, B, A);
//: interface  /sz:(225, 114) /bd:[ Ti0>A(36/225) Ti1>B(166/225) Ri0>Cin(52/114) Lo0<Cout(58/114) Bo0<S(117/225) ]
input B;    //: /sn:0 {0}(143,173)(159,173){1}
//: {2}(163,173)(176,173)(176,104)(186,104){3}
//: {4}(161,175)(161,176)(242,176)(242,152)(252,152){5}
input A;    //: /sn:0 {0}(130,98)(150,98){1}
//: {2}(154,98)(176,98)(176,99)(186,99){3}
//: {4}(152,100)(152,147)(252,147){5}
input Cin;    //: /sn:0 {0}(143,199)(213,199)(213,125){1}
//: {2}(215,123)(225,123)(225,124)(253,124){3}
//: {4}(213,121)(213,107)(223,107){5}
output Cout;    //: /sn:0 /dp:1 {0}(324,137)(347,137)(347,136)(357,136){1}
output S;    //: /sn:0 /dp:1 {0}(244,105)(348,105){1}
wire w4;    //: /sn:0 {0}(274,127)(293,127)(293,134)(303,134){1}
wire w2;    //: /sn:0 {0}(207,102)(215,102){1}
//: {2}(219,102)(223,102){3}
//: {4}(217,104)(217,129)(253,129){5}
wire w5;    //: /sn:0 {0}(273,150)(293,150)(293,139)(303,139){1}
//: enddecls

  //: output g4 (Cout) @(354,136) /sn:0 /w:[ 1 ]
  //: joint g8 (Cin) @(213, 123) /w:[ 2 4 -1 1 ]
  //: output g3 (S) @(345,105) /sn:0 /w:[ 1 ]
  //: input g2 (Cin) @(141,199) /sn:0 /w:[ 0 ]
  //: input g1 (B) @(141,173) /sn:0 /w:[ 0 ]
  and g10 (.I0(A), .I1(B), .Z(w5));   //: @(263,150) /sn:0 /tech:unit /w:[ 5 5 0 ]
  xor g6 (.I0(w2), .I1(Cin), .Z(S));   //: @(234,105) /sn:0 /delay:" 2" /w:[ 3 5 0 ]
  and g7 (.I0(Cin), .I1(w2), .Z(w4));   //: @(264,127) /sn:0 /tech:unit /w:[ 3 5 0 ]
  //: joint g9 (w2) @(217, 102) /w:[ 2 -1 1 4 ]
  //: joint g12 (B) @(161, 173) /w:[ 2 -1 1 4 ]
  xor g5 (.I0(A), .I1(B), .Z(w2));   //: @(197,102) /sn:0 /delay:" 2" /w:[ 3 3 0 ]
  //: joint g11 (A) @(152, 98) /w:[ 2 -1 1 4 ]
  //: input g0 (A) @(128,98) /sn:0 /w:[ 0 ]
  or g13 (.I0(w4), .I1(w5), .Z(Cout));   //: @(314,137) /sn:0 /tech:unit /w:[ 1 1 0 ]

endmodule

module main;    //: root_module
wire w13;    //: /sn:0 {0}(215,276)(215,266){1}
wire w6;    //: /sn:0 {0}(180,118)(180,128){1}
wire w7;    //: /sn:0 {0}(169,117)(169,128){1}
wire w4;    //: /sn:0 {0}(202,118)(202,128){1}
wire w3;    //: /sn:0 {0}(242,118)(242,128){1}
wire w0;    //: /sn:0 {0}(271,118)(271,128){1}
wire w12;    //: /sn:0 {0}(225,276)(225,266){1}
wire w10;    //: /sn:0 {0}(247,276)(247,266){1}
wire w1;    //: /sn:0 {0}(262,118)(262,128){1}
wire w8;    //: /sn:0 {0}(271,276)(271,266){1}
wire w14;    //: /sn:0 {0}(206,276)(206,266){1}
wire w11;    //: /sn:0 {0}(236,276)(236,266){1}
wire w2;    //: /sn:0 {0}(253,118)(253,128){1}
wire w15;    //: /sn:0 {0}(196,276)(196,266){1}
wire w5;    //: /sn:0 {0}(189,118)(189,128){1}
wire w9;    //: /sn:0 {0}(259,276)(259,266){1}
//: enddecls

  RCA_4b g0 (.Y3(w7), .Y2(w6), .Y1(w5), .Y0(w4), .X3(w3), .X2(w2), .X1(w1), .X0(w0), .Z7(w15), .Z6(w14), .Z5(w13), .Z4(w12), .Z3(w11), .Z2(w10), .Z1(w9), .Z0(w8));   //: @(155, 129) /sz:(128, 136) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Ti3>1 Ti4>1 Ti5>1 Ti6>1 Ti7>1 Bo0<1 Bo1<1 Bo2<1 Bo3<1 Bo4<1 Bo5<1 Bo6<1 Bo7<1 ]

endmodule
