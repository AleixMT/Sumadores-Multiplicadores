//: version "1.8.7"

module CarryLookahead_Logic(C2, P0, G0, P3, GG, G1, PG, P1, C3, Cout, P2, C1, G3, Cin, G2);
//: interface  /sz:(639, 96) /bd:[ Ti0>G0(557/639) Ti1>P0(520/639) Ti2>G1(409/639) Ti3>P1(368/639) Ti4>G2(270/639) Ti5>P2(227/639) Ti6>G3(107/639) Ti7>P3(54/639) Ri0>Cin(46/96) To0<C3(167/639) To1<C2(309/639) To2<C1(444/639) Lo0<Cout(39/96) Bo0<GG(545/639) Bo1<PG(472/639) ]
input G2;    //: /sn:0 {0}(370,94)(370,89){1}
//: {2}(372,87)(391,87)(391,405){3}
//: {4}(393,407)(653,407){5}
//: {6}(391,409)(391,517){7}
//: {8}(393,519)(553,519){9}
//: {10}(391,521)(391,739)(567,739){11}
//: {12}(370,85)(370,76)(371,76)(371,69){13}
output GG;    //: /sn:0 /dp:1 {0}(692,765)(708,765)(708,763)(718,763){1}
input P1;    //: /sn:0 {0}(569,809)(259,809)(259,686){1}
//: {2}(261,684)(564,684){3}
//: {4}(257,684)(255,684)(255,627){5}
//: {6}(257,625)(560,625){7}
//: {8}(255,623)(255,584){9}
//: {10}(257,582)(555,582){11}
//: {12}(255,580)(255,447)(245,447){13}
//: {14}(243,445)(243,422){15}
//: {16}(245,420)(549,420){17}
//: {18}(243,418)(243,325)(233,325){19}
//: {20}(231,323)(231,293){21}
//: {22}(233,291)(537,291){23}
//: {24}(231,289)(231,73){25}
//: {26}(231,327)(231,330)(543,330){27}
//: {28}(243,449)(243,450)(552,450){29}
output C3;    //: /sn:0 /dp:1 {0}(674,409)(712,409)(712,405)(722,405){1}
output PG;    //: /sn:0 /dp:1 {0}(585,681)(671,681){1}
input G0;    //: /sn:0 {0}(569,814)(205,814)(205,589){1}
//: {2}(207,587)(555,587){3}
//: {4}(205,585)(205,422)(195,422){5}
//: {6}(193,420)(193,298){7}
//: {8}(195,296)(537,296){9}
//: {10}(193,294)(193,199){11}
//: {12}(195,197)(540,197){13}
//: {14}(193,195)(193,70){15}
//: {16}(193,424)(193,425)(549,425){17}
output C2;    //: /sn:0 /dp:1 {0}(634,311)(642,311)(642,312)(652,312){1}
input Cin;    //: /sn:0 {0}(560,635)(83,635)(83,462){1}
//: {2}(85,460)(552,460){3}
//: {4}(83,458)(83,342){5}
//: {6}(85,340)(543,340){7}
//: {8}(83,338)(83,215){9}
//: {10}(85,213)(596,213){11}
//: {12}(83,211)(83,68){13}
input P3;    //: /sn:0 /dp:1 {0}(553,524)(433,524){1}
//: {2}(431,522)(431,64){3}
//: {4}(431,526)(431,542){5}
//: {6}(433,544)(556,544){7}
//: {8}(431,546)(431,570){9}
//: {10}(433,572)(555,572){11}
//: {12}(431,574)(431,613){13}
//: {14}(433,615)(560,615){15}
//: {16}(431,617)(431,672){17}
//: {18}(433,674)(564,674){19}
//: {20}(431,676)(431,732){21}
//: {22}(433,734)(567,734){23}
//: {24}(431,736)(431,765){25}
//: {26}(433,767)(569,767){27}
//: {28}(431,769)(431,799)(569,799){29}
input G1;    //: /sn:0 /dp:1 {0}(569,777)(279,777)(279,556){1}
//: {2}(281,554)(556,554){3}
//: {4}(279,552)(279,389){5}
//: {6}(281,387)(548,387){7}
//: {8}(279,385)(279,313){9}
//: {10}(281,311)(613,311){11}
//: {12}(279,309)(279,72){13}
output Cout;    //: /sn:0 /dp:1 {0}(686,553)(707,553)(707,545)(717,545){1}
input G3;    //: /sn:0 {0}(665,563)(492,563){1}
//: {2}(490,561)(490,63){3}
//: {4}(490,565)(490,763)(671,763){5}
output C1;    //: /sn:0 /dp:1 {0}(617,211)(626,211)(626,212)(636,212){1}
input P0;    //: /sn:0 {0}(564,689)(140,689)(140,632){1}
//: {2}(142,630)(560,630){3}
//: {4}(140,628)(140,457){5}
//: {6}(142,455)(552,455){7}
//: {8}(140,453)(140,337){9}
//: {10}(142,335)(543,335){11}
//: {12}(140,333)(140,204){13}
//: {14}(142,202)(540,202){15}
//: {16}(140,200)(140,69){17}
input P2;    //: /sn:0 /dp:1 {0}(548,382)(323,382){1}
//: {2}(321,380)(321,68){3}
//: {4}(321,384)(321,413){5}
//: {6}(323,415)(549,415){7}
//: {8}(321,417)(321,443){9}
//: {10}(323,445)(552,445){11}
//: {12}(321,447)(321,543){13}
//: {14}(319,545)(317,545)(317,575){15}
//: {16}(319,577)(555,577){17}
//: {18}(317,579)(317,618){19}
//: {20}(319,620)(560,620){21}
//: {22}(317,622)(317,674){23}
//: {24}(319,676)(329,676)(329,804)(569,804){25}
//: {26}(315,676)(305,676)(305,772)(569,772){27}
//: {28}(317,678)(317,679)(564,679){29}
//: {30}(321,547)(321,549)(556,549){31}
wire w6;    //: /sn:0 {0}(613,316)(574,316)(574,335)(564,335){1}
wire w4;    //: /sn:0 {0}(577,549)(620,549)(620,548)(665,548){1}
wire w3;    //: /sn:0 {0}(569,385)(643,385)(643,402)(653,402){1}
wire w0;    //: /sn:0 /dp:1 {0}(613,306)(568,306)(568,294)(558,294){1}
wire w12;    //: /sn:0 {0}(671,768)(600,768)(600,772)(590,772){1}
wire w1;    //: /sn:0 /dp:1 {0}(671,758)(598,758)(598,737)(588,737){1}
wire w8;    //: /sn:0 {0}(570,420)(643,420)(643,412)(653,412){1}
wire w17;    //: /sn:0 {0}(574,522)(655,522)(655,543)(665,543){1}
wire w14;    //: /sn:0 {0}(581,625)(642,625)(642,558)(665,558){1}
wire w11;    //: /sn:0 {0}(573,452)(650,452)(650,417)(653,417){1}
wire w15;    //: /sn:0 {0}(671,773)(618,773)(618,806)(590,806){1}
wire w5;    //: /sn:0 {0}(561,200)(586,200)(586,208)(596,208){1}
wire w9;    //: /sn:0 {0}(665,553)(633,553)(633,579)(576,579){1}
//: enddecls

  and g8 (.I0(P1), .I1(G0), .Z(w0));   //: @(548,294) /sn:0 /tech:unit /w:[ 23 9 1 ]
  or g4 (.I0(G0), .I1(P0), .Z(w5));   //: @(551,200) /sn:0 /tech:unit /w:[ 13 15 0 ]
  //: joint g44 (P1) @(243, 447) /w:[ 13 14 -1 28 ]
  or g16 (.I0(w0), .I1(G1), .I2(w6), .Z(C2));   //: @(624,311) /sn:0 /tech:unit /w:[ 0 11 0 0 ]
  and g3 (.I0(w5), .I1(Cin), .Z(C1));   //: @(607,211) /sn:0 /tech:unit /w:[ 1 11 0 ]
  //: joint g47 (P2) @(317, 577) /w:[ 16 15 -1 18 ]
  //: joint g26 (G0) @(193, 296) /w:[ 8 10 -1 7 ]
  //: output g17 (C2) @(649,312) /sn:0 /w:[ 1 ]
  //: input g2 (P0) @(140,67) /sn:0 /R:3 /w:[ 17 ]
  //: joint g30 (Cin) @(83, 340) /w:[ 6 8 -1 5 ]
  //: joint g23 (G1) @(279, 311) /w:[ 10 12 -1 9 ]
  //: joint g24 (P2) @(321, 382) /w:[ 1 2 -1 4 ]
  //: input g1 (G0) @(193,68) /sn:0 /R:3 /w:[ 15 ]
  //: joint g39 (P3) @(431, 524) /w:[ 1 2 -1 4 ]
  and g60 (.I0(P3), .I1(P2), .I2(G1), .Z(w12));   //: @(580,772) /sn:0 /w:[ 27 27 0 1 ]
  //: joint g29 (P0) @(140, 335) /w:[ 10 12 -1 9 ]
  or g51 (.I0(w17), .I1(w4), .I2(w9), .I3(w14), .I4(G3), .Z(Cout));   //: @(676,553) /sn:0 /w:[ 1 1 0 1 0 0 ]
  or g70 (.I0(w1), .I1(G3), .I2(w12), .I3(w15), .Z(GG));   //: @(682,765) /sn:0 /w:[ 0 5 0 0 0 ]
  //: input g18 (P3) @(431,62) /sn:0 /R:3 /w:[ 3 ]
  //: joint g65 (P1) @(259, 684) /w:[ 2 -1 4 1 ]
  //: joint g25 (P1) @(231, 325) /w:[ 19 20 -1 26 ]
  and g10 (.I0(P1), .I1(P0), .I2(Cin), .Z(w6));   //: @(554,335) /sn:0 /tech:unit /w:[ 27 11 7 1 ]
  //: joint g64 (P3) @(431, 734) /w:[ 22 21 -1 24 ]
  //: output g72 (GG) @(715,763) /sn:0 /w:[ 1 ]
  //: joint g49 (P0) @(140, 455) /w:[ 6 8 -1 5 ]
  //: input g6 (G1) @(279,70) /sn:0 /R:3 /w:[ 13 ]
  //: joint g50 (Cin) @(83, 460) /w:[ 2 4 -1 1 ]
  //: joint g68 (P2) @(317, 676) /w:[ 24 23 26 28 ]
  //: output g58 (PG) @(668,681) /sn:0 /w:[ 1 ]
  //: joint g56 (P1) @(255, 625) /w:[ 6 8 -1 5 ]
  and g35 (.I0(P3), .I1(P2), .I2(P1), .I3(G0), .Z(w9));   //: @(566,579) /sn:0 /w:[ 11 17 11 3 1 ]
  //: joint g9 (G0) @(193, 197) /w:[ 12 14 -1 11 ]
  //: input g7 (P1) @(231,71) /sn:0 /R:3 /w:[ 25 ]
  //: joint g71 (G3) @(490, 563) /w:[ 1 2 -1 4 ]
  and g59 (.I0(P3), .I1(G2), .Z(w1));   //: @(578,737) /sn:0 /w:[ 23 11 1 ]
  or g31 (.I0(w3), .I1(G2), .I2(w8), .I3(w11), .Z(C3));   //: @(664,409) /sn:0 /w:[ 1 5 1 1 0 ]
  and g22 (.I0(P2), .I1(P1), .I2(P0), .I3(Cin), .Z(w11));   //: @(563,452) /sn:0 /w:[ 11 29 7 3 0 ]
  //: joint g67 (P3) @(431, 767) /w:[ 26 25 -1 28 ]
  //: joint g54 (P3) @(431, 615) /w:[ 14 13 -1 16 ]
  and g36 (.I0(P3), .I1(P2), .I2(P1), .I3(P0), .I4(Cin), .Z(w14));   //: @(571,625) /sn:0 /w:[ 15 21 7 3 0 0 ]
  //: output g33 (C3) @(719,405) /sn:0 /w:[ 1 ]
  //: joint g41 (G1) @(279, 387) /w:[ 6 8 -1 5 ]
  //: joint g45 (G0) @(193, 422) /w:[ 5 6 -1 16 ]
  //: joint g69 (G0) @(205, 587) /w:[ 2 4 -1 1 ]
  //: joint g40 (P2) @(321, 445) /w:[ 10 9 -1 12 ]
  //: joint g42 (P3) @(431, 544) /w:[ 6 5 -1 8 ]
  //: output g52 (Cout) @(714,545) /sn:0 /w:[ 1 ]
  //: joint g66 (G1) @(279, 554) /w:[ 2 4 -1 1 ]
  //: input g12 (P2) @(321,66) /sn:0 /R:3 /w:[ 3 ]
  //: joint g57 (P0) @(140, 630) /w:[ 2 4 -1 1 ]
  and g34 (.I0(P3), .I1(P2), .I2(G1), .Z(w4));   //: @(567,549) /sn:0 /w:[ 7 31 3 0 ]
  //: joint g28 (P1) @(243, 420) /w:[ 16 18 -1 15 ]
  //: joint g46 (P3) @(431, 572) /w:[ 10 9 -1 12 ]
  //: joint g14 (P0) @(140, 202) /w:[ 14 16 -1 13 ]
  //: joint g11 (Cin) @(83, 213) /w:[ 10 12 -1 9 ]
  //: output g5 (C1) @(633,212) /sn:0 /w:[ 1 ]
  and g61 (.I0(P3), .I1(P2), .I2(P1), .I3(G0), .Z(w15));   //: @(580,806) /sn:0 /w:[ 29 25 0 0 1 ]
  and g21 (.I0(P2), .I1(P1), .I2(G0), .Z(w8));   //: @(560,420) /sn:0 /w:[ 7 17 17 0 ]
  //: input g19 (G3) @(490,61) /sn:0 /R:3 /w:[ 3 ]
  //: joint g32 (G2) @(370, 87) /w:[ 2 12 -1 1 ]
  and g20 (.I0(P2), .I1(G1), .Z(w3));   //: @(559,385) /sn:0 /w:[ 0 7 0 ]
  //: joint g63 (G2) @(391, 519) /w:[ 8 7 -1 10 ]
  //: joint g38 (G2) @(391, 407) /w:[ 4 3 -1 6 ]
  //: joint g15 (P1) @(231, 291) /w:[ 22 24 -1 21 ]
  //: input g0 (Cin) @(83,66) /sn:0 /R:3 /w:[ 13 ]
  //: joint g43 (P2) @(321, 545) /w:[ -1 13 14 30 ]
  //: joint g27 (P2) @(321, 415) /w:[ 6 5 -1 8 ]
  //: joint g48 (P1) @(255, 582) /w:[ 10 12 -1 9 ]
  //: joint g62 (P3) @(431, 674) /w:[ 18 17 -1 20 ]
  and g37 (.I0(G2), .I1(P3), .Z(w17));   //: @(564,522) /sn:0 /w:[ 9 0 0 ]
  //: joint g55 (P2) @(317, 620) /w:[ 20 19 -1 22 ]
  and g53 (.I0(P3), .I1(P2), .I2(P1), .I3(P0), .Z(PG));   //: @(575,681) /sn:0 /w:[ 19 29 3 0 0 ]
  //: input g13 (G2) @(371,67) /sn:0 /R:3 /w:[ 13 ]

endmodule

module CLA_Adder_4bit(S0, A1, S3, A0, A2, B1, S1, P, A3, S2, Cin, B0, B2, G, B3);
//: interface  /sz:(209, 138) /bd:[ Ti0>B3(42/209) Ti1>B2(63/209) Ti2>B1(79/209) Ti3>B0(99/209) Ti4>A3(130/209) Ti5>A2(151/209) Ti6>A1(172/209) Ti7>A0(190/209) Bi0>S3(14/209) Bi1>S2(38/209) Ri0>Cin(59/138) Bo0<S1(61/209) Bo1<S0(87/209) Bo2<G(148/209) Bo3<P(119/209) ]
input A0;    //: /sn:0 {0}(986,200)(986,255)(990,255)(990,272){1}
output S1;    //: /sn:0 /dp:1 {0}(808,460)(808,450)(809,450)(809,391){1}
input A3;    //: /sn:0 {0}(419,190)(462,190)(462,265){1}
output G;    //: /sn:0 {0}(887,612)(887,656){1}
input A2;    //: /sn:0 {0}(629,177)(629,252)(631,252)(631,274){1}
input B2;    //: /sn:0 {0}(579,183)(579,267)(580,267)(580,274){1}
input Cin;    //: /sn:0 {0}(1187,305)(1077,305)(1077,325){1}
//: {2}(1075,327)(1034,327)(1034,329)(1028,329){3}
//: {4}(1077,329)(1077,561)(982,561){5}
input B1;    //: /sn:0 {0}(766,208)(766,274){1}
output S0;    //: /sn:0 /dp:1 {0}(1000,520)(1000,389){1}
output P;    //: /sn:0 {0}(814,612)(814,660){1}
input A1;    //: /sn:0 {0}(809,198)(809,274){1}
input B3;    //: /sn:0 {0}(348,220)(406,220)(406,265){1}
output S3;    //: /sn:0 {0}(462,458)(462,382){1}
input B0;    //: /sn:0 {0}(898,176)(931,176)(931,272){1}
output S2;    //: /sn:0 /dp:1 {0}(647,459)(647,435)(635,435)(635,391){1}
wire w16;    //: /sn:0 /dp:1 {0}(569,514)(569,506)(547,506)(547,391){1}
wire w34;    //: /sn:0 /dp:1 {0}(663,331)(684,331)(684,486)(651,486)(651,514){1}
wire w4;    //: /sn:0 /dp:1 {0}(862,514)(862,441)(919,441)(919,389){1}
wire w22;    //: /sn:0 /dp:1 {0}(396,514)(396,506)(374,506)(374,382){1}
wire w3;    //: /sn:0 /dp:1 {0}(899,514)(899,506)(957,506)(957,389){1}
wire w10;    //: /sn:0 /dp:1 {0}(710,514)(710,474)(721,474)(721,391){1}
wire w21;    //: /sn:0 /dp:1 {0}(449,514)(449,506)(419,506)(419,382){1}
wire w33;    //: /sn:0 {0}(786,514)(786,479)(855,479)(855,331)(837,331){1}
wire w35;    //: /sn:0 {0}(509,514)(509,322)(490,322){1}
wire w2;    //: /sn:0 {0}(341,554)(308,554)(308,494){1}
wire w15;    //: /sn:0 /dp:1 {0}(612,514)(612,488)(592,488)(592,391){1}
wire w9;    //: /sn:0 /dp:1 {0}(751,514)(751,434)(766,434)(766,391){1}
//: enddecls

  CarryLookahead_Logic g4 (.G0(w3), .P0(w4), .G1(w9), .P1(w10), .G2(w15), .P2(w16), .G3(w21), .P3(w22), .Cin(Cin), .C3(w35), .C2(w34), .C1(w33), .Cout(w2), .GG(G), .PG(P));   //: @(342, 515) /sz:(639, 96) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>0 Ti3>0 Ti4>0 Ti5>0 Ti6>0 Ti7>0 Ri0>5 To0<0 To1<1 To2<0 Lo0<0 Bo0<0 Bo1<0 ]
  //: output g44 (S0) @(1000,517) /sn:0 /R:3 /w:[ 0 ]
  //: input g8 (A1) @(809,196) /sn:0 /R:3 /w:[ 0 ]
  PFA_v1 g3 (.A(A3), .B(B3), .C(w35), .S(S3), .P(w22), .G(w21));   //: @(363, 266) /sz:(126, 115) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Bo0<1 Bo1<1 Bo2<1 ]
  //: output g47 (S3) @(462,455) /sn:0 /R:3 /w:[ 0 ]
  //: input g16 (A0) @(986,198) /sn:0 /R:3 /w:[ 0 ]
  PFA_v1 g2 (.A(A2), .B(B2), .C(w34), .S(S2), .P(w16), .G(w15));   //: @(536, 275) /sz:(126, 115) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Bo0<1 Bo1<1 Bo2<1 ]
  PFA_v1 g1 (.A(A1), .B(B1), .C(w33), .S(S1), .P(w10), .G(w9));   //: @(710, 275) /sz:(126, 115) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Bo0<1 Bo1<1 Bo2<1 ]
  //: input g10 (A2) @(629,175) /sn:0 /R:3 /w:[ 0 ]
  //: joint g6 (Cin) @(1077, 327) /w:[ -1 1 2 4 ]
  led g7 (.I(w2));   //: @(308,487) /sn:0 /w:[ 1 ] /type:0
  //: input g9 (B1) @(766,206) /sn:0 /R:3 /w:[ 0 ]
  //: output g45 (S1) @(808,457) /sn:0 /R:3 /w:[ 0 ]
  //: output g42 (P) @(814,657) /sn:0 /R:3 /w:[ 1 ]
  //: input g12 (A3) @(417,190) /sn:0 /w:[ 0 ]
  //: output g46 (S2) @(647,456) /sn:0 /R:3 /w:[ 0 ]
  //: input g5 (Cin) @(1189,305) /sn:0 /R:2 /w:[ 0 ]
  //: input g14 (B0) @(896,176) /sn:0 /w:[ 0 ]
  //: input g11 (B2) @(579,181) /sn:0 /R:3 /w:[ 0 ]
  PFA_v1 g0 (.A(A0), .B(B0), .C(Cin), .S(S0), .P(w4), .G(w3));   //: @(901, 273) /sz:(126, 115) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>3 Bo0<1 Bo1<1 Bo2<1 ]
  //: output g43 (G) @(887,653) /sn:0 /R:3 /w:[ 1 ]
  //: input g13 (B3) @(346,220) /sn:0 /w:[ 0 ]

endmodule

module PFA_v1(C, B, P, S, A, G);
//: interface  /sz:(126, 115) /bd:[ Ti0>A(21/126) Ti1>B(82/126) Ri0>C(56/115) Bo0<S(99/126) Bo1<P(11/126) Bo2<G(56/126) ]
input B;    //: /sn:0 {0}(144,200)(161,200){1}
//: {2}(165,200)(202,200)(202,177)(210,177){3}
//: {4}(163,202)(163,320){5}
//: {6}(165,322)(231,322){7}
//: {8}(163,324)(163,361)(240,361){9}
input A;    //: /sn:0 {0}(151,147)(178,147){1}
//: {2}(182,147)(202,147)(202,172)(210,172){3}
//: {4}(180,149)(180,317)(188,317){5}
//: {6}(192,317)(231,317){7}
//: {8}(190,319)(190,356)(240,356){9}
output G;    //: /sn:0 /dp:1 {0}(261,359)(337,359)(337,385)(346,385){1}
input C;    //: /sn:0 {0}(149,271)(266,271)(266,186)(276,186){1}
output P;    //: /sn:0 /dp:1 {0}(252,320)(312,320)(312,319)(322,319){1}
output S;    //: /sn:0 /dp:1 {0}(297,184)(394,184)(394,198)(406,198){1}
wire w2;    //: /sn:0 {0}(231,175)(267,175)(267,181)(276,181){1}
//: enddecls

  xor g4 (.I0(w2), .I1(C), .Z(S));   //: @(287,184) /sn:0 /delay:" 2" /w:[ 1 1 0 ]
  //: joint g8 (B) @(163, 200) /w:[ 2 -1 1 4 ]
  xor g3 (.I0(A), .I1(B), .Z(w2));   //: @(221,175) /sn:0 /delay:" 2" /w:[ 3 3 0 ]
  //: input g2 (C) @(147,271) /sn:0 /w:[ 0 ]
  //: input g1 (B) @(142,200) /sn:0 /w:[ 0 ]
  and g10 (.I0(A), .I1(B), .Z(G));   //: @(251,359) /sn:0 /delay:" 1" /w:[ 9 9 0 ]
  or g6 (.I0(A), .I1(B), .Z(P));   //: @(242,320) /sn:0 /delay:" 1" /w:[ 7 7 0 ]
  //: joint g7 (A) @(180, 147) /w:[ 2 -1 1 4 ]
  //: output g9 (P) @(319,319) /sn:0 /w:[ 1 ]
  //: joint g12 (A) @(190, 317) /w:[ 6 -1 5 8 ]
  //: output g5 (S) @(403,198) /sn:0 /w:[ 1 ]
  //: joint g11 (B) @(163, 322) /w:[ 6 5 -1 8 ]
  //: input g0 (A) @(149,147) /sn:0 /w:[ 0 ]
  //: output g13 (G) @(343,385) /sn:0 /w:[ 1 ]

endmodule

module main;    //: root_module
wire w16;    //: /sn:0 /dp:1 {0}(-93,687)(-93,618)(6,618)(6,522){1}
wire w58;    //: /sn:0 {0}(84,785)(84,813)(101,813)(101,817){1}
wire w65;    //: /sn:0 {0}(-345,164)(-270,164)(-270,391){1}
wire w50;    //: /sn:0 {0}(-55,159)(17,159)(17,398){1}
wire w59;    //: /sn:0 {0}(-86,292)(-71,292)(-71,398){1}
wire w81;    //: /sn:0 {0}(-52,522)(-52,826)(-76,826)(-76,913){1}
wire w25;    //: /sn:0 {0}(236,123)(356,123)(356,366){1}
wire w62;    //: /sn:0 {0}(-345,135)(-249,135)(-249,391){1}
wire w72;    //: /sn:0 {0}(-662,196)(-601,196)(-601,381){1}
wire w39;    //: /sn:0 {0}(-75,522)(-75,809)(-133,809)(-133,906){1}
wire w3;    //: /sn:0 {0}(271,506)(271,876)(170,876)(170,910){1}
wire w0;    //: /sn:0 {0}(245,506)(245,868)(118,868)(118,909){1}
wire w36;    //: /sn:0 {0}(-386,531)(-386,928)(-384,928)(-384,941){1}
wire w60;    //: /sn:0 {0}(-86,259)(-50,259)(-50,398){1}
wire w20;    //: /sn:0 {0}(-495,899)(-495,784)(-639,784)(-639,521){1}
wire w30;    //: /sn:0 {0}(303,506)(303,641)(59,641)(59,687){1}
wire w29;    //: /sn:0 {0}(237,153)(335,153)(335,366){1}
wire w71;    //: /sn:0 {0}(-634,103)(-528,103)(-528,381){1}
wire w66;    //: /sn:0 {0}(-375,233)(-321,233)(-321,391){1}
wire w73;    //: /sn:0 {0}(-633,162)(-570,162)(-570,381){1}
wire w63;    //: /sn:0 {0}(-346,105)(-228,105)(-228,391){1}
wire w54;    //: /sn:0 {0}(-152,687)(-152,451)(-190,451){1}
wire w70;    //: /sn:0 {0}(-633,133)(-549,133)(-549,381){1}
wire w31;    //: /sn:0 {0}(332,506)(332,664)(96,664)(96,687){1}
wire w1;    //: /sn:0 {0}(222,506)(222,863)(56,863)(56,908){1}
wire w68;    //: /sn:0 {0}(-376,264)(-337,264)(-337,391){1}
wire w32;    //: /sn:0 {0}(-662,521)(-662,798)(-552,798)(-552,892){1}
wire w53;    //: /sn:0 {0}(-17,687)(-17,684)(55,684)(55,591)(166,591)(166,451)(97,451){1}
wire w46;    //: /sn:0 {0}(207,251)(263,251)(263,366){1}
wire w8;    //: /sn:0 {0}(-503,713)(-503,727)(-462,727){1}
wire w52;    //: /sn:0 {0}(179,734)(456,734)(456,425){1}
//: {2}(458,423)(489,423)(489,433)(497,433){3}
//: {4}(454,423)(428,423)(428,426)(394,426){5}
wire w44;    //: /sn:0 {0}(208,216)(283,216)(283,366){1}
wire w27;    //: /sn:0 {0}(-57,70)(77,70)(77,398){1}
wire w75;    //: /sn:0 {0}(-664,295)(-658,295)(-658,381){1}
wire w28;    //: /sn:0 {0}(-56,100)(59,100)(59,398){1}
wire w67;    //: /sn:0 {0}(-376,297)(-358,297)(-358,391){1}
wire w80;    //: /sn:0 {0}(-26,522)(-26,835)(-24,835)(-24,914){1}
wire w35;    //: /sn:0 {0}(-362,531)(-362,852)(-336,852)(-336,932){1}
wire w14;    //: /sn:0 {0}(235,93)(374,93)(374,366){1}
wire w45;    //: /sn:0 {0}(206,282)(247,282)(247,366){1}
wire w49;    //: /sn:0 {0}(-84,193)(-14,193)(-14,398){1}
wire w69;    //: /sn:0 {0}(-635,73)(-510,73)(-510,381){1}
wire w41;    //: /sn:0 {0}(237,182)(314,182)(314,366){1}
wire w48;    //: /sn:0 {0}(-55,130)(38,130)(38,398){1}
wire w74;    //: /sn:0 {0}(-663,231)(-621,231)(-621,381){1}
wire w2;    //: /sn:0 {0}(198,506)(198,856)(13,856)(13,911){1}
wire w78;    //: /sn:0 {0}(-313,531)(-313,827)(-227,827)(-227,940){1}
wire w47;    //: /sn:0 {0}(206,315)(226,315)(226,366){1}
wire w15;    //: /sn:0 /dp:1 {0}(-52,687)(-52,650)(35,650)(35,522){1}
wire w85;    //: /sn:0 {0}(-613,521)(-613,772)(-443,772)(-443,900){1}
wire w55;    //: /sn:0 {0}(-317,687)(-317,629)(-449,629)(-449,441)(-490,441){1}
wire w61;    //: /sn:0 {0}(-347,75)(-210,75)(-210,391){1}
wire w38;    //: /sn:0 {0}(-686,521)(-686,814)(-600,814)(-600,901){1}
wire w64;    //: /sn:0 {0}(-374,198)(-301,198)(-301,391){1}
wire w87;    //: /sn:0 /dp:1 {0}(-407,687)(-407,605)(-581,605)(-581,521){1}
wire w43;    //: /sn:0 /dp:1 {0}(-354,687)(-354,657)(-367,657)(-367,645)(-552,645)(-552,521){1}
wire w76;    //: /sn:0 {0}(-664,262)(-637,262)(-637,381){1}
wire w26;    //: /sn:0 /dp:1 {0}(-234,687)(-234,568)(-281,568)(-281,531){1}
wire w57;    //: /sn:0 {0}(11,785)(11,816)(21,816)(21,820){1}
wire w51;    //: /sn:0 {0}(-85,228)(-34,228)(-34,398){1}
wire w40;    //: /sn:0 {0}(-99,522)(-99,797)(-181,797)(-181,915){1}
wire w77;    //: /sn:0 {0}(-252,531)(-252,550)(-191,550)(-191,687){1}
wire w79;    //: /sn:0 {0}(-339,531)(-339,843)(-279,843)(-279,939){1}
//: enddecls

  led g4 (.I(w58));   //: @(101,824) /sn:0 /R:2 /w:[ 1 ] /type:0
  //: switch g8 (w14) @(218,93) /sn:0 /w:[ 0 ] /st:0
  led g44 (.I(w36));   //: @(-384,948) /sn:0 /R:2 /w:[ 1 ] /type:0
  CarryLookahead_Logic g3 (.G0(w31), .P0(w30), .G1(w15), .P1(w16), .G2(w77), .P2(w26), .G3(w43), .P3(w87), .Cin(w52), .C3(w55), .C2(w54), .C1(w53), .Cout(w8), .GG(w58), .PG(w57));   //: @(-461, 688) /sz:(639, 96) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>0 Ti3>0 Ti4>1 Ti5>0 Ti6>0 Ti7>0 Ri0>0 To0<0 To1<0 To2<0 Lo0<1 Bo0<0 Bo1<0 ]
  //: switch g16 (w27) @(-74,70) /sn:0 /w:[ 0 ] /st:0
  led g47 (.I(w81));   //: @(-76,920) /sn:0 /R:2 /w:[ 1 ] /type:0
  //: switch g17 (w48) @(-72,130) /sn:0 /w:[ 0 ] /st:0
  //: switch g26 (w63) @(-363,105) /sn:0 /w:[ 0 ] /st:0
  led g2 (.I(w1));   //: @(56,915) /sn:0 /R:2 /w:[ 1 ] /type:0
  //: switch g23 (w60) @(-103,259) /sn:0 /w:[ 0 ] /st:0
  //: switch g30 (w67) @(-393,297) /sn:0 /w:[ 0 ] /st:0
  //: switch g24 (w61) @(-364,75) /sn:0 /w:[ 0 ] /st:0
  //: switch g39 (w76) @(-681,262) /sn:0 /w:[ 0 ] /st:0
  led g1 (.I(w0));   //: @(118,916) /sn:0 /R:2 /w:[ 1 ] /type:0
  //: switch g29 (w66) @(-392,233) /sn:0 /w:[ 0 ] /st:0
  led g51 (.I(w20));   //: @(-495,906) /sn:0 /R:2 /w:[ 0 ] /type:0
  //: switch g18 (w28) @(-73,100) /sn:0 /w:[ 0 ] /st:0
  //: switch g10 (w29) @(220,153) /sn:0 /w:[ 0 ] /st:0
  //: switch g25 (w62) @(-362,135) /sn:0 /w:[ 0 ] /st:0
  led g49 (.I(w80));   //: @(-24,921) /sn:0 /R:2 /w:[ 1 ] /type:0
  //: switch g6 (w52) @(515,433) /sn:0 /R:2 /w:[ 3 ] /st:0
  led g50 (.I(w32));   //: @(-552,899) /sn:0 /R:2 /w:[ 1 ] /type:0
  //: joint g7 (w52) @(456, 423) /w:[ 2 -1 4 1 ]
  //: switch g9 (w25) @(219,123) /sn:0 /w:[ 0 ] /st:0
  //: switch g35 (w72) @(-679,196) /sn:0 /w:[ 0 ] /st:0
  CLA_Adder_4bit g56 (.B3(w75), .B2(w76), .B1(w74), .B0(w72), .A3(w73), .A2(w70), .A1(w71), .A0(w69), .S3(w38), .S2(w32), .Cin(w55), .S1(w20), .S0(w85), .G(w43), .P(w87));   //: @(-700, 382) /sz:(209, 138) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Ti3>1 Ti4>1 Ti5>1 Ti6>1 Ti7>1 Bi0>0 Bi1>0 Ri0>1 Bo0<1 Bo1<0 Bo2<1 Bo3<1 ]
  //: switch g22 (w59) @(-103,292) /sn:0 /w:[ 0 ] /st:0
  //: switch g31 (w68) @(-393,264) /sn:0 /w:[ 0 ] /st:0
  //: switch g33 (w70) @(-650,133) /sn:0 /w:[ 0 ] /st:0
  //: switch g36 (w73) @(-650,162) /sn:0 /w:[ 0 ] /st:0
  led g41 (.I(w35));   //: @(-336,939) /sn:0 /R:2 /w:[ 1 ] /type:0
  led g45 (.I(w78));   //: @(-227,947) /sn:0 /R:2 /w:[ 1 ] /type:0
  CLA_Adder_4bit g54 (.B3(w59), .B2(w60), .B1(w51), .B0(w49), .A3(w50), .A2(w48), .A1(w28), .A0(w27), .S3(w40), .S2(w39), .Cin(w53), .S1(w81), .S0(w80), .G(w15), .P(w16));   //: @(-113, 399) /sz:(209, 122) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Ti3>1 Ti4>1 Ti5>1 Ti6>1 Ti7>1 Bi0>0 Bi1>0 Ri0>1 Bo0<0 Bo1<0 Bo2<1 Bo3<1 ]
  CLA_Adder_4bit g42 (.B3(w47), .B2(w45), .B1(w46), .B0(w44), .A3(w41), .A2(w29), .A1(w25), .A0(w14), .S3(w2), .S2(w1), .Cin(w52), .S1(w0), .S0(w3), .G(w31), .P(w30));   //: @(184, 367) /sz:(209, 138) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Ti3>1 Ti4>1 Ti5>1 Ti6>1 Ti7>1 Bi0>0 Bi1>0 Ri0>5 Bo0<0 Bo1<0 Bo2<0 Bo3<0 ]
  led g40 (.I(w2));   //: @(13,918) /sn:0 /R:2 /w:[ 1 ] /type:0
  led g52 (.I(w38));   //: @(-600,908) /sn:0 /R:2 /w:[ 1 ] /type:0
  //: switch g12 (w44) @(191,216) /sn:0 /w:[ 0 ] /st:0
  //: switch g28 (w65) @(-362,164) /sn:0 /w:[ 0 ] /st:0
  //: switch g34 (w71) @(-651,103) /sn:0 /w:[ 0 ] /st:0
  led g46 (.I(w39));   //: @(-133,913) /sn:0 /R:2 /w:[ 1 ] /type:0
  led g57 (.I(w8));   //: @(-503,706) /sn:0 /w:[ 0 ] /type:0
  led g5 (.I(w57));   //: @(21,827) /sn:0 /R:2 /w:[ 1 ] /type:0
  //: switch g11 (w41) @(220,182) /sn:0 /w:[ 0 ] /st:0
  //: switch g14 (w46) @(190,251) /sn:0 /w:[ 0 ] /st:0
  //: switch g19 (w49) @(-101,193) /sn:0 /w:[ 0 ] /st:0
  //: switch g21 (w51) @(-102,228) /sn:0 /w:[ 0 ] /st:0
  //: switch g20 (w50) @(-72,159) /sn:0 /w:[ 0 ] /st:0
  //: switch g32 (w69) @(-652,73) /sn:0 /w:[ 0 ] /st:0
  //: switch g15 (w47) @(189,315) /sn:0 /w:[ 0 ] /st:0
  //: switch g38 (w75) @(-681,295) /sn:0 /w:[ 0 ] /st:0
  led g0 (.I(w3));   //: @(170,917) /sn:0 /R:2 /w:[ 1 ] /type:0
  led g43 (.I(w79));   //: @(-279,946) /sn:0 /R:2 /w:[ 1 ] /type:0
  //: switch g27 (w64) @(-391,198) /sn:0 /w:[ 0 ] /st:0
  led g48 (.I(w40));   //: @(-181,922) /sn:0 /R:2 /w:[ 1 ] /type:0
  //: switch g37 (w74) @(-680,231) /sn:0 /w:[ 0 ] /st:0
  CLA_Adder_4bit g55 (.B3(w67), .B2(w68), .B1(w66), .B0(w64), .A3(w65), .A2(w62), .A1(w63), .A0(w61), .S3(w36), .S2(w35), .Cin(w54), .S1(w79), .S0(w78), .G(w77), .P(w26));   //: @(-400, 392) /sz:(209, 138) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Ti3>1 Ti4>1 Ti5>1 Ti6>1 Ti7>1 Bi0>0 Bi1>0 Ri0>1 Bo0<0 Bo1<0 Bo2<0 Bo3<1 ]
  //: switch g13 (w45) @(189,282) /sn:0 /w:[ 0 ] /st:0
  led g53 (.I(w85));   //: @(-443,907) /sn:0 /R:2 /w:[ 1 ] /type:0

endmodule
