//: version "1.8.7"

module CarryLookahead_Logic(C2, P0, G0, P3, GG, G1, PG, P1, C3, Cout, P2, C1, G3, Cin, G2);
//: interface  /sz:(639, 96) /bd:[ Ti0>G0(557/639) Ti1>P0(520/639) Ti2>G1(409/639) Ti3>P1(368/639) Ti4>G2(270/639) Ti5>P2(227/639) Ti6>G3(107/639) Ti7>P3(54/639) Ri0>Cin(46/96) To0<C3(167/639) To1<C2(309/639) To2<C1(444/639) Lo0<Cout(39/96) Bo0<GG(545/639) Bo1<PG(472/639) ]
input G2;    //: /sn:0 {0}(370,94)(370,89){1}
//: {2}(372,87)(391,87)(391,405){3}
//: {4}(393,407)(653,407){5}
//: {6}(391,409)(391,517){7}
//: {8}(393,519)(553,519){9}
//: {10}(391,521)(391,739)(567,739){11}
//: {12}(370,85)(370,76)(371,76)(371,69){13}
output GG;    //: /sn:0 /dp:1 {0}(692,761)(708,761)(708,763)(718,763){1}
input P1;    //: /sn:0 {0}(569,809)(259,809)(259,686){1}
//: {2}(261,684)(564,684){3}
//: {4}(257,684)(255,684)(255,627){5}
//: {6}(257,625)(560,625){7}
//: {8}(255,623)(255,584){9}
//: {10}(257,582)(555,582){11}
//: {12}(255,580)(255,447)(245,447){13}
//: {14}(243,445)(243,422){15}
//: {16}(245,420)(549,420){17}
//: {18}(243,418)(243,325)(233,325){19}
//: {20}(231,323)(231,293){21}
//: {22}(233,291)(537,291){23}
//: {24}(231,289)(231,73){25}
//: {26}(231,327)(231,330)(544,330){27}
//: {28}(243,449)(243,450)(552,450){29}
output C3;    //: /sn:0 /dp:1 {0}(674,409)(712,409)(712,405)(722,405){1}
output PG;    //: /sn:0 /dp:1 {0}(585,681)(671,681){1}
input G0;    //: /sn:0 {0}(569,814)(205,814)(205,589){1}
//: {2}(207,587)(555,587){3}
//: {4}(205,585)(205,422)(195,422){5}
//: {6}(193,420)(193,298){7}
//: {8}(195,296)(537,296){9}
//: {10}(193,294)(193,199){11}
//: {12}(193,195)(193,70){13}
//: {14}(191,197)(180,197)(180,194)(537,194){15}
//: {16}(193,424)(193,425)(549,425){17}
output C2;    //: /sn:0 /dp:1 {0}(634,311)(642,311)(642,312)(652,312){1}
input Cin;    //: /sn:0 {0}(560,635)(83,635)(83,462){1}
//: {2}(85,460)(552,460){3}
//: {4}(83,458)(83,342){5}
//: {6}(85,340)(544,340){7}
//: {8}(83,338)(83,215){9}
//: {10}(83,211)(83,68){11}
//: {12}(81,213)(72,213)(72,214)(585,214){13}
input P3;    //: /sn:0 /dp:1 {0}(553,524)(433,524){1}
//: {2}(431,522)(431,64){3}
//: {4}(431,526)(431,542){5}
//: {6}(433,544)(556,544){7}
//: {8}(431,546)(431,570){9}
//: {10}(433,572)(555,572){11}
//: {12}(431,574)(431,613){13}
//: {14}(433,615)(560,615){15}
//: {16}(431,617)(431,672){17}
//: {18}(433,674)(564,674){19}
//: {20}(431,676)(431,732){21}
//: {22}(433,734)(567,734){23}
//: {24}(431,736)(431,765){25}
//: {26}(433,767)(569,767){27}
//: {28}(431,769)(431,799)(569,799){29}
input G1;    //: /sn:0 /dp:1 {0}(569,777)(279,777)(279,556){1}
//: {2}(281,554)(556,554){3}
//: {4}(279,552)(279,389){5}
//: {6}(281,387)(548,387){7}
//: {8}(279,385)(279,313){9}
//: {10}(281,311)(613,311){11}
//: {12}(279,309)(279,72){13}
output Cout;    //: /sn:0 /dp:1 {0}(688,554)(709,554)(709,545)(717,545){1}
input G3;    //: /sn:0 {0}(667,564)(580,564)(580,563)(492,563){1}
//: {2}(490,561)(490,63){3}
//: {4}(490,565)(490,759)(671,759){5}
output C1;    //: /sn:0 /dp:1 {0}(606,212)(636,212){1}
input P0;    //: /sn:0 {0}(564,689)(140,689)(140,632){1}
//: {2}(142,630)(560,630){3}
//: {4}(140,628)(140,457){5}
//: {6}(142,455)(552,455){7}
//: {8}(140,453)(140,337){9}
//: {10}(142,335)(544,335){11}
//: {12}(140,333)(140,204){13}
//: {14}(142,202)(153,202)(153,189)(358,189)(358,199)(537,199){15}
//: {16}(140,200)(140,69){17}
input P2;    //: /sn:0 /dp:1 {0}(548,382)(323,382){1}
//: {2}(321,380)(321,68){3}
//: {4}(321,384)(321,413){5}
//: {6}(323,415)(549,415){7}
//: {8}(321,417)(321,443){9}
//: {10}(323,445)(552,445){11}
//: {12}(321,447)(321,543){13}
//: {14}(319,545)(317,545)(317,575){15}
//: {16}(319,577)(555,577){17}
//: {18}(317,579)(317,618){19}
//: {20}(319,620)(560,620){21}
//: {22}(317,622)(317,674){23}
//: {24}(319,676)(329,676)(329,804)(569,804){25}
//: {26}(315,676)(305,676)(305,772)(569,772){27}
//: {28}(317,678)(317,679)(564,679){29}
//: {30}(321,547)(321,549)(556,549){31}
wire w6;    //: /sn:0 {0}(613,316)(575,316)(575,335)(565,335){1}
wire w4;    //: /sn:0 {0}(577,549)(667,549){1}
wire w3;    //: /sn:0 {0}(569,385)(643,385)(643,402)(653,402){1}
wire w0;    //: /sn:0 /dp:1 {0}(613,306)(568,306)(568,294)(558,294){1}
wire w12;    //: /sn:0 {0}(671,764)(600,764)(600,772)(590,772){1}
wire w10;    //: /sn:0 {0}(558,197)(574,197)(574,209)(585,209){1}
wire w1;    //: /sn:0 /dp:1 {0}(671,754)(598,754)(598,737)(588,737){1}
wire w8;    //: /sn:0 {0}(570,420)(643,420)(643,412)(653,412){1}
wire w17;    //: /sn:0 {0}(574,522)(657,522)(657,544)(667,544){1}
wire w14;    //: /sn:0 {0}(581,625)(644,625)(644,559)(667,559){1}
wire w11;    //: /sn:0 {0}(573,452)(650,452)(650,417)(653,417){1}
wire w15;    //: /sn:0 {0}(671,769)(618,769)(618,806)(590,806){1}
wire w9;    //: /sn:0 {0}(667,554)(635,554)(635,579)(576,579){1}
//: enddecls

  or g4 (.I0(w10), .I1(Cin), .Z(C1));   //: @(596,212) /sn:0 /tech:unit /w:[ 1 13 0 ]
  and g8 (.I0(P1), .I1(G0), .Z(w0));   //: @(548,294) /sn:0 /tech:unit /w:[ 23 9 1 ]
  //: joint g44 (P1) @(243, 447) /w:[ 13 14 -1 28 ]
  or g16 (.I0(w0), .I1(G1), .I2(w6), .Z(C2));   //: @(624,311) /sn:0 /tech:unit /w:[ 0 11 0 0 ]
  //: joint g47 (P2) @(317, 577) /w:[ 16 15 -1 18 ]
  //: joint g26 (G0) @(193, 296) /w:[ 8 10 -1 7 ]
  //: output g17 (C2) @(649,312) /sn:0 /w:[ 1 ]
  //: input g2 (P0) @(140,67) /sn:0 /R:3 /w:[ 17 ]
  //: joint g30 (Cin) @(83, 340) /w:[ 6 8 -1 5 ]
  //: joint g23 (G1) @(279, 311) /w:[ 10 12 -1 9 ]
  //: joint g24 (P2) @(321, 382) /w:[ 1 2 -1 4 ]
  //: input g1 (G0) @(193,68) /sn:0 /R:3 /w:[ 13 ]
  //: joint g39 (P3) @(431, 524) /w:[ 1 2 -1 4 ]
  and g60 (.I0(P3), .I1(P2), .I2(G1), .Z(w12));   //: @(580,772) /sn:0 /tech:unit /w:[ 27 27 0 1 ]
  //: joint g29 (P0) @(140, 335) /w:[ 10 12 -1 9 ]
  or g51 (.I0(w17), .I1(w4), .I2(w9), .I3(w14), .I4(G3), .Z(Cout));   //: @(678,554) /sn:0 /tech:unit /w:[ 1 1 0 1 0 0 ]
  or g70 (.I0(w1), .I1(G3), .I2(w12), .I3(w15), .Z(GG));   //: @(682,761) /sn:0 /tech:unit /w:[ 0 5 0 0 0 ]
  //: input g18 (P3) @(431,62) /sn:0 /R:3 /w:[ 3 ]
  //: joint g65 (P1) @(259, 684) /w:[ 2 -1 4 1 ]
  //: joint g25 (P1) @(231, 325) /w:[ 19 20 -1 26 ]
  and g10 (.I0(P1), .I1(P0), .I2(Cin), .Z(w6));   //: @(555,335) /sn:0 /tech:unit /w:[ 27 11 7 1 ]
  //: joint g64 (P3) @(431, 734) /w:[ 22 21 -1 24 ]
  //: output g72 (GG) @(715,763) /sn:0 /w:[ 1 ]
  //: joint g49 (P0) @(140, 455) /w:[ 6 8 -1 5 ]
  //: input g6 (G1) @(279,70) /sn:0 /R:3 /w:[ 13 ]
  //: joint g50 (Cin) @(83, 460) /w:[ 2 4 -1 1 ]
  and g73 (.I0(G0), .I1(P0), .Z(w10));   //: @(548,197) /sn:0 /tech:unit /w:[ 15 15 0 ]
  //: joint g68 (P2) @(317, 676) /w:[ 24 23 26 28 ]
  //: output g58 (PG) @(668,681) /sn:0 /w:[ 1 ]
  //: joint g56 (P1) @(255, 625) /w:[ 6 8 -1 5 ]
  and g35 (.I0(P3), .I1(P2), .I2(P1), .I3(G0), .Z(w9));   //: @(566,579) /sn:0 /tech:unit /w:[ 11 17 11 3 1 ]
  //: joint g9 (G0) @(193, 197) /w:[ -1 12 14 11 ]
  //: input g7 (P1) @(231,71) /sn:0 /R:3 /w:[ 25 ]
  //: joint g71 (G3) @(490, 563) /w:[ 1 2 -1 4 ]
  and g59 (.I0(P3), .I1(G2), .Z(w1));   //: @(578,737) /sn:0 /tech:unit /w:[ 23 11 1 ]
  or g31 (.I0(w3), .I1(G2), .I2(w8), .I3(w11), .Z(C3));   //: @(664,409) /sn:0 /tech:unit /w:[ 1 5 1 1 0 ]
  and g22 (.I0(P2), .I1(P1), .I2(P0), .I3(Cin), .Z(w11));   //: @(563,452) /sn:0 /tech:unit /w:[ 11 29 7 3 0 ]
  //: joint g67 (P3) @(431, 767) /w:[ 26 25 -1 28 ]
  //: joint g54 (P3) @(431, 615) /w:[ 14 13 -1 16 ]
  and g36 (.I0(P3), .I1(P2), .I2(P1), .I3(P0), .I4(Cin), .Z(w14));   //: @(571,625) /sn:0 /tech:unit /w:[ 15 21 7 3 0 0 ]
  //: output g33 (C3) @(719,405) /sn:0 /w:[ 1 ]
  //: joint g41 (G1) @(279, 387) /w:[ 6 8 -1 5 ]
  //: joint g45 (G0) @(193, 422) /w:[ 5 6 -1 16 ]
  //: joint g69 (G0) @(205, 587) /w:[ 2 4 -1 1 ]
  //: joint g40 (P2) @(321, 445) /w:[ 10 9 -1 12 ]
  //: joint g42 (P3) @(431, 544) /w:[ 6 5 -1 8 ]
  //: output g52 (Cout) @(714,545) /sn:0 /w:[ 1 ]
  //: joint g66 (G1) @(279, 554) /w:[ 2 4 -1 1 ]
  //: input g12 (P2) @(321,66) /sn:0 /R:3 /w:[ 3 ]
  //: joint g57 (P0) @(140, 630) /w:[ 2 4 -1 1 ]
  and g34 (.I0(P3), .I1(P2), .I2(G1), .Z(w4));   //: @(567,549) /sn:0 /tech:unit /w:[ 7 31 3 0 ]
  //: joint g28 (P1) @(243, 420) /w:[ 16 18 -1 15 ]
  //: joint g46 (P3) @(431, 572) /w:[ 10 9 -1 12 ]
  //: joint g14 (P0) @(140, 202) /w:[ 14 16 -1 13 ]
  //: joint g11 (Cin) @(83, 213) /w:[ -1 10 12 9 ]
  //: output g5 (C1) @(633,212) /sn:0 /w:[ 1 ]
  and g61 (.I0(P3), .I1(P2), .I2(P1), .I3(G0), .Z(w15));   //: @(580,806) /sn:0 /tech:unit /w:[ 29 25 0 0 1 ]
  and g21 (.I0(P2), .I1(P1), .I2(G0), .Z(w8));   //: @(560,420) /sn:0 /tech:unit /w:[ 7 17 17 0 ]
  //: input g19 (G3) @(490,61) /sn:0 /R:3 /w:[ 3 ]
  //: joint g32 (G2) @(370, 87) /w:[ 2 12 -1 1 ]
  and g20 (.I0(P2), .I1(G1), .Z(w3));   //: @(559,385) /sn:0 /tech:unit /w:[ 0 7 0 ]
  //: joint g63 (G2) @(391, 519) /w:[ 8 7 -1 10 ]
  //: joint g38 (G2) @(391, 407) /w:[ 4 3 -1 6 ]
  //: joint g15 (P1) @(231, 291) /w:[ 22 24 -1 21 ]
  //: input g0 (Cin) @(83,66) /sn:0 /R:3 /w:[ 11 ]
  //: joint g43 (P2) @(321, 545) /w:[ -1 13 14 30 ]
  //: joint g27 (P2) @(321, 415) /w:[ 6 5 -1 8 ]
  //: joint g48 (P1) @(255, 582) /w:[ 10 12 -1 9 ]
  //: joint g62 (P3) @(431, 674) /w:[ 18 17 -1 20 ]
  and g37 (.I0(G2), .I1(P3), .Z(w17));   //: @(564,522) /sn:0 /tech:unit /w:[ 9 0 0 ]
  //: joint g55 (P2) @(317, 620) /w:[ 20 19 -1 22 ]
  and g53 (.I0(P3), .I1(P2), .I2(P1), .I3(P0), .Z(PG));   //: @(575,681) /sn:0 /tech:unit /w:[ 19 29 3 0 0 ]
  //: input g13 (G2) @(371,67) /sn:0 /R:3 /w:[ 13 ]

endmodule

module CLA_Adder_4bit(S0, A1, S3, A0, A2, B1, S1, P, A3, S2, Cin, B0, B2, G, B3);
//: interface  /sz:(209, 138) /bd:[ Ti0>B3(42/209) Ti1>B2(63/209) Ti2>B1(79/209) Ti3>B0(99/209) Ti4>A3(130/209) Ti5>A2(151/209) Ti6>A1(172/209) Ti7>A0(190/209) Bi0>S3(14/209) Bi1>S2(38/209) Ri0>Cin(59/138) Bo0<S1(61/209) Bo1<S0(87/209) Bo2<G(148/209) Bo3<P(119/209) ]
input A0;    //: /sn:0 {0}(986,200)(986,235){1}
//: {2}(988,237)(1003,237)(1003,224){3}
//: {4}(986,239)(986,257)(990,257)(990,272){5}
output S1;    //: /sn:0 /dp:1 {0}(808,460)(808,452)(809,452)(809,428){1}
//: {2}(809,424)(809,391){3}
//: {4}(807,426)(790,426)(790,419){5}
input A3;    //: /sn:0 {0}(419,190)(462,190)(462,230){1}
//: {2}(464,232)(471,232)(471,222){3}
//: {4}(462,234)(462,265){5}
output G;    //: /sn:0 {0}(887,612)(887,632){1}
//: {2}(889,634)(909,634)(909,632){3}
//: {4}(887,636)(887,656){5}
input A2;    //: /sn:0 {0}(629,177)(629,215){1}
//: {2}(631,217)(652,217)(652,206){3}
//: {4}(629,219)(629,254)(631,254)(631,274){5}
input B2;    //: /sn:0 {0}(579,183)(579,223){1}
//: {2}(581,225)(596,225)(596,214){3}
//: {4}(579,227)(579,269)(580,269)(580,274){5}
input Cin;    //: /sn:0 {0}(1187,305)(1077,305)(1077,325){1}
//: {2}(1075,327)(1034,327)(1034,329)(1028,329){3}
//: {4}(1077,329)(1077,521){5}
//: {6}(1079,523)(1106,523)(1106,510){7}
//: {8}(1077,525)(1077,561)(982,561){9}
input B1;    //: /sn:0 {0}(766,208)(766,228){1}
//: {2}(768,230)(788,230)(788,212){3}
//: {4}(766,232)(766,274){5}
output S0;    //: /sn:0 /dp:1 {0}(1000,520)(1000,457){1}
//: {2}(1002,455)(1018,455)(1018,447){3}
//: {4}(1000,453)(1000,389){5}
output P;    //: /sn:0 {0}(814,612)(814,639){1}
//: {2}(816,641)(842,641)(842,631){3}
//: {4}(814,643)(814,660){5}
input A1;    //: /sn:0 {0}(809,198)(809,241){1}
//: {2}(811,243)(833,243)(833,233){3}
//: {4}(809,245)(809,274){5}
input B3;    //: /sn:0 {0}(348,220)(406,220)(406,245){1}
//: {2}(408,247)(424,247)(424,236){3}
//: {4}(406,249)(406,265){5}
output S3;    //: /sn:0 {0}(462,458)(462,435){1}
//: {2}(462,431)(462,382){3}
//: {4}(460,433)(448,433)(448,422){5}
input B0;    //: /sn:0 {0}(898,176)(931,176)(931,245){1}
//: {2}(933,247)(948,247)(948,228){3}
//: {4}(931,249)(931,272){5}
output S2;    //: /sn:0 /dp:1 {0}(647,459)(647,437)(635,437)(635,432){1}
//: {2}(635,428)(635,391){3}
//: {4}(633,430)(605,430)(605,423){5}
wire w16;    //: /sn:0 /dp:1 {0}(569,514)(569,508)(547,508)(547,473){1}
//: {2}(547,469)(547,391){3}
//: {4}(545,471)(527,471)(527,455){5}
wire w34;    //: /sn:0 /dp:1 {0}(663,331)(684,331)(684,452){1}
//: {2}(682,454)(670,454)(670,446){3}
//: {4}(684,456)(684,488)(651,488)(651,514){5}
wire w4;    //: /sn:0 /dp:1 {0}(862,514)(862,481){1}
//: {2}(864,479)(905,479)(905,469){3}
//: {4}(862,477)(862,439)(919,439)(919,389){5}
wire w22;    //: /sn:0 /dp:1 {0}(396,514)(396,508)(374,508)(374,424){1}
//: {2}(374,420)(374,382){3}
//: {4}(372,422)(341,422)(341,411){5}
wire w3;    //: /sn:0 /dp:1 {0}(899,514)(899,508)(957,508)(957,473){1}
//: {2}(959,471)(967,471)(967,454){3}
//: {4}(957,469)(957,389){5}
wire w10;    //: /sn:0 /dp:1 {0}(710,514)(710,476)(721,476)(721,438){1}
//: {2}(721,434)(721,391){3}
//: {4}(719,436)(694,436)(694,429){5}
wire w21;    //: /sn:0 /dp:1 {0}(449,514)(449,508)(419,508)(419,451){1}
//: {2}(419,447)(419,382){3}
//: {4}(417,449)(398,449)(398,438){5}
wire w33;    //: /sn:0 {0}(786,514)(786,481)(855,481)(855,423){1}
//: {2}(857,421)(868,421)(868,415){3}
//: {4}(855,419)(855,331)(837,331){5}
wire w35;    //: /sn:0 {0}(509,514)(509,443){1}
//: {2}(509,439)(509,322)(490,322){3}
//: {4}(507,441)(489,441)(489,428){5}
wire w2;    //: /sn:0 {0}(341,554)(308,554)(308,494){1}
wire w15;    //: /sn:0 /dp:1 {0}(612,514)(612,490)(592,490)(592,451){1}
//: {2}(592,447)(592,391){3}
//: {4}(590,449)(578,449)(578,461)(563,461)(563,451){5}
wire w9;    //: /sn:0 /dp:1 {0}(751,514)(751,463){1}
//: {2}(751,459)(751,432)(766,432)(766,391){3}
//: {4}(749,461)(733,461)(733,452){5}
//: enddecls

  CarryLookahead_Logic g4 (.G0(w3), .P0(w4), .G1(w9), .P1(w10), .G2(w15), .P2(w16), .G3(w21), .P3(w22), .Cin(Cin), .C3(w35), .C2(w34), .C1(w33), .Cout(w2), .GG(G), .PG(P));   //: @(342, 515) /sz:(639, 96) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>0 Ti3>0 Ti4>0 Ti5>0 Ti6>0 Ti7>0 Ri0>9 To0<0 To1<5 To2<0 Lo0<0 Bo0<0 Bo1<0 ]
  //: output g44 (S0) @(1000,517) /sn:0 /R:3 /w:[ 0 ]
  //: input g8 (A1) @(809,196) /sn:0 /R:3 /w:[ 0 ]
  PFA_v1 g3 (.A(A3), .B(B3), .C(w35), .S(S3), .P(w22), .G(w21));   //: @(363, 266) /sz:(126, 115) /sn:0 /p:[ Ti0>5 Ti1>5 Ri0>3 Bo0<3 Bo1<3 Bo2<3 ]
  //: output g47 (S3) @(462,455) /sn:0 /R:3 /w:[ 0 ]
  //: input g16 (A0) @(986,198) /sn:0 /R:3 /w:[ 0 ]
  //: joint g17 (S0) @(1000, 455) /w:[ 2 4 -1 1 ]
  led g26 (.I(w9));   //: @(733,445) /sn:0 /w:[ 5 ] /type:0
  PFA_v1 g2 (.A(A2), .B(B2), .C(w34), .S(S2), .P(w16), .G(w15));   //: @(536, 275) /sz:(126, 115) /sn:0 /p:[ Ti0>5 Ti1>5 Ri0>0 Bo0<3 Bo1<3 Bo2<3 ]
  //: joint g23 (w33) @(855, 421) /w:[ 2 4 -1 1 ]
  led g30 (.I(w34));   //: @(670,439) /sn:0 /w:[ 3 ] /type:0
  PFA_v1 g1 (.A(A1), .B(B1), .C(w33), .S(S1), .P(w10), .G(w9));   //: @(710, 275) /sz:(126, 115) /sn:0 /p:[ Ti0>5 Ti1>5 Ri0>5 Bo0<3 Bo1<3 Bo2<3 ]
  led g24 (.I(S1));   //: @(790,412) /sn:0 /w:[ 5 ] /type:0
  //: joint g39 (w35) @(509, 441) /w:[ -1 2 4 1 ]
  //: joint g29 (w10) @(721, 436) /w:[ -1 2 4 1 ]
  led g60 (.I(B0));   //: @(948,221) /sn:0 /w:[ 3 ] /type:0
  //: joint g51 (w22) @(374, 422) /w:[ -1 2 4 1 ]
  led g18 (.I(w3));   //: @(967,447) /sn:0 /w:[ 3 ] /type:0
  led g70 (.I(A3));   //: @(471,215) /sn:0 /w:[ 3 ] /type:0
  //: input g10 (A2) @(629,175) /sn:0 /R:3 /w:[ 0 ]
  //: joint g25 (S1) @(809, 426) /w:[ -1 2 4 1 ]
  //: joint g65 (B1) @(766, 230) /w:[ 2 1 -1 4 ]
  led g64 (.I(B1));   //: @(788,205) /sn:0 /w:[ 3 ] /type:0
  //: joint g49 (w21) @(419, 449) /w:[ -1 2 4 1 ]
  led g72 (.I(B3));   //: @(424,229) /sn:0 /w:[ 3 ] /type:0
  //: joint g6 (Cin) @(1077, 327) /w:[ -1 1 2 4 ]
  led g50 (.I(w22));   //: @(341,404) /sn:0 /w:[ 5 ] /type:0
  led g7 (.I(w2));   //: @(308,487) /sn:0 /w:[ 1 ] /type:0
  //: input g9 (B1) @(766,206) /sn:0 /R:3 /w:[ 0 ]
  //: joint g35 (w15) @(592, 449) /w:[ -1 2 4 1 ]
  led g56 (.I(Cin));   //: @(1106,503) /sn:0 /w:[ 7 ] /type:0
  led g58 (.I(A0));   //: @(1003,217) /sn:0 /w:[ 3 ] /type:0
  led g68 (.I(B2));   //: @(596,207) /sn:0 /w:[ 3 ] /type:0
  //: joint g73 (B3) @(406, 247) /w:[ 2 1 -1 4 ]
  led g22 (.I(w33));   //: @(868,408) /sn:0 /w:[ 3 ] /type:0
  //: joint g31 (w34) @(684, 454) /w:[ -1 1 2 4 ]
  //: joint g59 (A0) @(986, 237) /w:[ 2 1 -1 4 ]
  //: joint g71 (A3) @(462, 232) /w:[ 2 1 -1 4 ]
  //: joint g67 (A2) @(629, 217) /w:[ 2 1 -1 4 ]
  //: output g45 (S1) @(808,457) /sn:0 /R:3 /w:[ 0 ]
  //: joint g33 (S2) @(635, 430) /w:[ -1 2 4 1 ]
  led g36 (.I(w16));   //: @(527,448) /sn:0 /w:[ 5 ] /type:0
  //: joint g41 (S3) @(462, 433) /w:[ -1 2 4 1 ]
  led g54 (.I(G));   //: @(909,625) /sn:0 /w:[ 3 ] /type:0
  //: output g42 (P) @(814,657) /sn:0 /R:3 /w:[ 5 ]
  led g40 (.I(S3));   //: @(448,415) /sn:0 /w:[ 5 ] /type:0
  led g52 (.I(P));   //: @(842,624) /sn:0 /w:[ 3 ] /type:0
  //: joint g69 (B2) @(579, 225) /w:[ 2 1 -1 4 ]
  led g66 (.I(A2));   //: @(652,199) /sn:0 /w:[ 3 ] /type:0
  //: input g12 (A3) @(417,190) /sn:0 /w:[ 0 ]
  //: output g46 (S2) @(647,456) /sn:0 /R:3 /w:[ 0 ]
  led g28 (.I(w10));   //: @(694,422) /sn:0 /w:[ 5 ] /type:0
  led g34 (.I(w15));   //: @(563,444) /sn:0 /w:[ 5 ] /type:0
  //: joint g57 (Cin) @(1077, 523) /w:[ 6 5 -1 8 ]
  //: input g5 (Cin) @(1189,305) /sn:0 /R:2 /w:[ 0 ]
  //: input g14 (B0) @(896,176) /sn:0 /w:[ 0 ]
  //: input g11 (B2) @(579,181) /sn:0 /R:3 /w:[ 0 ]
  //: joint g19 (w3) @(957, 471) /w:[ 2 4 -1 1 ]
  //: joint g21 (w4) @(862, 479) /w:[ 2 4 -1 1 ]
  //: joint g61 (B0) @(931, 247) /w:[ 2 1 -1 4 ]
  led g20 (.I(w4));   //: @(905,462) /sn:0 /w:[ 3 ] /type:0
  led g32 (.I(S2));   //: @(605,416) /sn:0 /w:[ 5 ] /type:0
  //: joint g63 (A1) @(809, 243) /w:[ 2 1 -1 4 ]
  PFA_v1 g0 (.A(A0), .B(B0), .C(Cin), .S(S0), .P(w4), .G(w3));   //: @(901, 273) /sz:(126, 115) /sn:0 /p:[ Ti0>5 Ti1>5 Ri0>3 Bo0<5 Bo1<5 Bo2<5 ]
  //: output g43 (G) @(887,653) /sn:0 /R:3 /w:[ 5 ]
  led g15 (.I(S0));   //: @(1018,440) /sn:0 /w:[ 3 ] /type:0
  led g38 (.I(w35));   //: @(489,421) /sn:0 /w:[ 5 ] /type:0
  //: joint g27 (w9) @(751, 461) /w:[ -1 2 4 1 ]
  led g48 (.I(w21));   //: @(398,431) /sn:0 /w:[ 5 ] /type:0
  //: joint g37 (w16) @(547, 471) /w:[ -1 2 4 1 ]
  led g62 (.I(A1));   //: @(833,226) /sn:0 /w:[ 3 ] /type:0
  //: joint g55 (G) @(887, 634) /w:[ 2 1 -1 4 ]
  //: input g13 (B3) @(346,220) /sn:0 /w:[ 0 ]
  //: joint g53 (P) @(814, 641) /w:[ 2 1 -1 4 ]

endmodule

module PFA_v1(C, B, P, S, A, G);
//: interface  /sz:(126, 115) /bd:[ Ti0>A(21/126) Ti1>B(82/126) Ri0>C(56/115) Bo0<S(99/126) Bo1<P(11/126) Bo2<G(56/126) ]
input B;    //: /sn:0 {0}(144,200)(161,200){1}
//: {2}(165,200)(202,200)(202,177)(210,177){3}
//: {4}(163,202)(163,320){5}
//: {6}(165,322)(231,322){7}
//: {8}(163,324)(163,361)(240,361){9}
input A;    //: /sn:0 {0}(151,147)(178,147){1}
//: {2}(182,147)(202,147)(202,172)(210,172){3}
//: {4}(180,149)(180,317)(188,317){5}
//: {6}(192,317)(231,317){7}
//: {8}(190,319)(190,356)(240,356){9}
output G;    //: /sn:0 /dp:1 {0}(261,359)(337,359)(337,385)(346,385){1}
input C;    //: /sn:0 {0}(149,271)(266,271)(266,186)(276,186){1}
output P;    //: /sn:0 /dp:1 {0}(252,320)(312,320)(312,319)(322,319){1}
output S;    //: /sn:0 /dp:1 {0}(297,184)(394,184)(394,198)(406,198){1}
wire w2;    //: /sn:0 {0}(231,175)(267,175)(267,181)(276,181){1}
//: enddecls

  xor g4 (.I0(w2), .I1(C), .Z(S));   //: @(287,184) /sn:0 /delay:" 2" /w:[ 1 1 0 ]
  //: joint g8 (B) @(163, 200) /w:[ 2 -1 1 4 ]
  xor g3 (.I0(A), .I1(B), .Z(w2));   //: @(221,175) /sn:0 /delay:" 2" /w:[ 3 3 0 ]
  //: input g2 (C) @(147,271) /sn:0 /w:[ 0 ]
  //: input g1 (B) @(142,200) /sn:0 /w:[ 0 ]
  and g10 (.I0(A), .I1(B), .Z(G));   //: @(251,359) /sn:0 /delay:" 1" /w:[ 9 9 0 ]
  or g6 (.I0(A), .I1(B), .Z(P));   //: @(242,320) /sn:0 /delay:" 1" /w:[ 7 7 0 ]
  //: joint g7 (A) @(180, 147) /w:[ 2 -1 1 4 ]
  //: output g9 (P) @(319,319) /sn:0 /w:[ 1 ]
  //: joint g12 (A) @(190, 317) /w:[ 6 -1 5 8 ]
  //: output g5 (S) @(403,198) /sn:0 /w:[ 1 ]
  //: joint g11 (B) @(163, 322) /w:[ 6 5 -1 8 ]
  //: input g0 (A) @(149,147) /sn:0 /w:[ 0 ]
  //: output g13 (G) @(343,385) /sn:0 /w:[ 1 ]

endmodule

module main;    //: root_module
wire w16;    //: /sn:0 {0}(1088,243)(1088,237)(1066,237)(1066,202){1}
//: {2}(1066,198)(1066,120){3}
//: {4}(1064,200)(1046,200)(1046,184){5}
wire w6;    //: /sn:0 {0}(590,468)(590,435){1}
//: {2}(592,433)(633,433)(633,423){3}
//: {4}(590,431)(590,393)(647,393)(647,343){5}
wire w13;    //: /sn:0 {0}(-205,683)(-205,650){1}
//: {2}(-203,648)(-162,648)(-162,638){3}
//: {4}(-205,646)(-205,608)(-148,608)(-148,558){5}
wire S1;    //: /sn:0 {0}(1309,148)(1309,155)(1328,155)(1328,120){1}
wire w7;    //: /sn:0 {0}(-978,841)(-978,835)(-920,835)(-920,800){1}
//: {2}(-918,798)(-910,798)(-910,781){3}
//: {4}(-920,796)(-920,716){5}
wire w58;    //: /sn:0 {0}(-1111,-109)(925,-109)(925,-26){1}
//: {2}(927,-24)(943,-24)(943,-35){3}
//: {4}(925,-22)(925,-6){5}
wire w65;    //: /sn:0 {0}(-1366,-216)(-626,-216)(-626,401)(-607,401){1}
//: {2}(-603,401)(-596,401)(-596,391){3}
//: {4}(-605,403)(-605,434){5}
wire w34;    //: /sn:0 {0}(1182,60)(1203,60)(1203,181){1}
//: {2}(1201,183)(1189,183)(1189,175){3}
//: {4}(1203,185)(1203,217)(1170,217)(1170,243){5}
wire G2;    //: /sn:0 {0}(-990,939)(-990,961)(-968,961)(-968,959){1}
wire w50;    //: /sn:0 {0}(-1394,10)(-682,10)(-682,419)(-663,419){1}
//: {2}(-661,417)(-661,414)(-643,414)(-643,405){3}
//: {4}(-661,421)(-661,434){5}
wire w59;    //: /sn:0 {0}(-1075,-123)(1085,-123)(1085,-39)(1096,-39){1}
//: {2}(1098,-41)(1098,-48)(1115,-48)(1115,-57){3}
//: {4}(1098,-37)(1098,0)(1099,0)(1099,3){5}
wire w4;    //: /sn:0 {0}(1381,243)(1381,210){1}
//: {2}(1383,208)(1424,208)(1424,198){3}
//: {4}(1381,206)(1381,168)(1438,168)(1438,118){5}
wire S6;    //: /sn:0 {0}(333,377)(333,384)(363,384)(363,345){1}
wire S7;    //: /sn:0 {0}(518,373)(518,380)(537,380)(537,345){1}
wire w25;    //: /sn:0 {0}(-498,683)(-498,677)(-520,677)(-520,642){1}
//: {2}(-520,638)(-520,560){3}
//: {4}(-522,640)(-540,640)(-540,624){5}
wire Cin1;    //: /sn:0 {0}(39,679)(39,692)(12,692){1}
//: {2}(10,690)(10,500){3}
//: {4}(12,498)(34,498){5}
//: {6}(36,496)(36,448){7}
//: {8}(36,500)(36,508)(69,508){9}
//: {10}(8,498)(-39,498){11}
//: {12}(10,694)(10,730)(-85,730){13}
wire w39;    //: /sn:0 {0}(-558,683)(-558,612){1}
//: {2}(-558,608)(-558,491)(-577,491){3}
//: {4}(-560,610)(-578,610)(-578,597){5}
wire P1;    //: /sn:0 {0}(-253,781)(-253,810)(-225,810)(-225,800){1}
wire w62;    //: /sn:0 {0}(-1403,-201)(-912,-201)(-912,564)(-893,564){1}
//: {2}(-889,564)(-874,564)(-874,551){3}
//: {4}(-891,566)(-891,586)(-887,586)(-887,599){5}
wire w72;    //: /sn:0 {0}(-1119,-320)(714,-320)(714,189){1}
//: {2}(716,191)(731,191)(731,178){3}
//: {4}(714,193)(714,213)(718,213)(718,226){5}
wire w56;    //: /sn:0 {0}(-1182,-79)(494,-79)(494,182){1}
//: {2}(496,184)(516,184)(516,166){3}
//: {4}(494,186)(494,228){5}
wire w3;    //: /sn:0 {0}(1418,243)(1418,237)(1476,237)(1476,202){1}
//: {2}(1478,200)(1486,200)(1486,183){3}
//: {4}(1476,198)(1476,118){5}
wire w22;    //: /sn:0 {0}(915,243)(915,237)(893,237)(893,153){1}
//: {2}(893,149)(893,111){3}
//: {4}(891,151)(860,151)(860,140){5}
wire w36;    //: /sn:0 {0}(237,468)(237,397){1}
//: {2}(237,393)(237,276)(218,276){3}
//: {4}(235,395)(217,395)(217,382){5}
wire w0;    //: /sn:0 {0}(1668,55)(1608,55)(1608,56)(1598,56){1}
//: {2}(1594,56)(1551,56)(1551,58)(1547,58){3}
//: {4}(1596,58)(1596,250){5}
//: {6}(1598,252)(1625,252)(1625,239){7}
//: {8}(1596,254)(1596,290)(1501,290){9}
wire w20;    //: /sn:0 {0}(-455,683)(-455,659)(-475,659)(-475,620){1}
//: {2}(-475,616)(-475,560){3}
//: {4}(-477,618)(-489,618)(-489,630)(-504,630)(-504,620){5}
wire w60;    //: /sn:0 {0}(-1040,-137)(1285,-137)(1285,-43){1}
//: {2}(1287,-41)(1307,-41)(1307,-59){3}
//: {4}(1285,-39)(1285,3){5}
wire w29;    //: /sn:0 {0}(-1126,841)(-1126,790){1}
//: {2}(-1126,786)(-1126,759)(-1111,759)(-1111,718){3}
//: {4}(-1128,788)(-1144,788)(-1144,779){5}
wire w30;    //: /sn:0 {0}(-1167,841)(-1167,803)(-1156,803)(-1156,765){1}
//: {2}(-1156,761)(-1156,718){3}
//: {4}(-1158,763)(-1183,763)(-1183,756){5}
wire w71;    //: /sn:0 {0}(-1296,-247)(-258,-247)(-258,410){1}
//: {2}(-256,412)(-234,412)(-234,402){3}
//: {4}(-258,414)(-258,443){5}
wire w37;    //: /sn:0 {0}(391,285)(412,285)(412,406){1}
//: {2}(410,408)(398,408)(398,400){3}
//: {4}(412,410)(412,442)(379,442)(379,468){5}
wire w42;    //: /sn:0 {0}(-1428,841)(-1428,835)(-1458,835)(-1458,778){1}
//: {2}(-1458,774)(-1458,709){3}
//: {4}(-1460,776)(-1479,776)(-1479,765){5}
wire Cin2;    //: /sn:0 {0}(-895,888)(-800,888)(-800,666){1}
//: {2}(-798,664)(-783,664)(-783,687)(-761,687){3}
//: {4}(-759,685)(-759,663){5}
//: {6}(-759,689)(-759,723)(-726,723){7}
//: {8}(-800,662)(-800,656)(-849,656){9}
wire G;    //: /sn:0 {0}(1406,341)(1406,363)(1428,363)(1428,361){1}
wire w12;    //: /sn:0 {0}(438,468)(438,430)(449,430)(449,392){1}
//: {2}(449,388)(449,345){3}
//: {4}(447,390)(422,390)(422,383){5}
wire w18;    //: /sn:0 {0}(297,468)(297,462)(275,462)(275,427){1}
//: {2}(275,423)(275,345){3}
//: {4}(273,425)(255,425)(255,409){5}
wire S4;    //: /sn:0 {0}(728,343)(728,409)(746,409)(746,401){1}
wire w19;    //: /sn:0 {0}(-357,683)(-357,645)(-346,645)(-346,607){1}
//: {2}(-346,603)(-346,560){3}
//: {4}(-348,605)(-373,605)(-373,598){5}
wire w66;    //: /sn:0 {0}(-1439,-184)(-1068,-184)(-1068,568){1}
//: {2}(-1066,570)(-1044,570)(-1044,560){3}
//: {4}(-1068,572)(-1068,601){5}
wire w73;    //: /sn:0 {0}(-1047,-349)(1135,-349)(1135,-54)(1146,-54){1}
//: {2}(1150,-54)(1171,-54)(1171,-65){3}
//: {4}(1148,-52)(1148,-15)(1150,-15)(1150,3){5}
wire w10;    //: /sn:0 {0}(1229,243)(1229,205)(1240,205)(1240,167){1}
//: {2}(1240,163)(1240,120){3}
//: {4}(1238,165)(1213,165)(1213,158){5}
wire w23;    //: /sn:0 {0}(177,468)(177,462)(147,462)(147,405){1}
//: {2}(147,401)(147,336){3}
//: {4}(145,403)(126,403)(126,392){5}
wire G0;    //: /sn:0 {0}(615,566)(615,588)(637,588)(637,586){1}
wire w63;    //: /sn:0 {0}(-1512,-154)(-1415,-154)(-1415,557){1}
//: {2}(-1413,559)(-1406,559)(-1406,549){3}
//: {4}(-1415,561)(-1415,592){5}
wire S8;    //: /sn:0 {0}(-67,558)(-67,624)(-49,624)(-49,616){1}
wire S9;    //: /sn:0 {0}(-619,591)(-619,602)(-605,602)(-605,551){1}
wire w54;    //: /sn:0 {0}(-1253,-49)(134,-49)(134,199){1}
//: {2}(136,201)(152,201)(152,190){3}
//: {4}(134,203)(134,219){5}
wire w70;    //: /sn:0 {0}(-1012,-363)(1328,-363)(1328,-30){1}
//: {2}(1330,-28)(1352,-28)(1352,-38){3}
//: {4}(1328,-26)(1328,3){5}
wire w21;    //: /sn:0 {0}(968,243)(968,237)(938,237)(938,180){1}
//: {2}(938,176)(938,111){3}
//: {4}(936,178)(917,178)(917,167){5}
wire w24;    //: /sn:0 {0}(124,468)(124,462)(102,462)(102,378){1}
//: {2}(102,374)(102,336){3}
//: {4}(100,376)(69,376)(69,365){5}
wire Cin0;    //: /sn:0 {0}(834,464)(834,477)(807,477){1}
//: {2}(805,475)(805,285){3}
//: {4}(807,283)(832,283)(832,281){5}
//: {6}(834,283)(860,283){7}
//: {8}(830,283)(827,283)(827,223){9}
//: {10}(803,283)(756,283){11}
//: {12}(805,479)(805,515)(710,515){13}
wire S11;    //: /sn:0 {0}(-277,588)(-277,595)(-258,595)(-258,560){1}
wire w31;    //: /sn:0 {0}(-1265,841)(-1265,817)(-1285,817)(-1285,778){1}
//: {2}(-1285,774)(-1285,718){3}
//: {4}(-1287,776)(-1299,776)(-1299,788)(-1314,788)(-1314,778){5}
wire w1;    //: /sn:0 {0}(-1540,72)(-1471,72)(-1471,572){1}
//: {2}(-1469,574)(-1453,574)(-1453,563){3}
//: {4}(-1471,576)(-1471,592){5}
wire S0;    //: /sn:0 {0}(1519,118)(1519,184)(1537,184)(1537,176){1}
wire w32;    //: /sn:0 {0}(-1308,841)(-1308,835)(-1330,835)(-1330,800){1}
//: {2}(-1330,796)(-1330,718){3}
//: {4}(-1332,798)(-1350,798)(-1350,782){5}
wire w68;    //: /sn:0 {0}(-1154,-305)(537,-305)(537,195){1}
//: {2}(539,197)(561,197)(561,187){3}
//: {4}(537,199)(537,228){5}
wire S5;    //: /sn:0 {0}(176,376)(176,387)(190,387)(190,336){1}
wire w53;    //: /sn:0 {0}(-1289,-35)(-136,-35)(-136,414){1}
//: {2}(-134,416)(-119,416)(-119,397){3}
//: {4}(-136,418)(-136,441){5}
wire w8;    //: /sn:0 {0}(-168,683)(-168,677)(-110,677)(-110,642){1}
//: {2}(-108,640)(-100,640)(-100,623){3}
//: {4}(-110,638)(-110,558){5}
wire w46;    //: /sn:0 {0}(-1091,841)(-1091,808)(-1022,808)(-1022,750){1}
//: {2}(-1020,748)(-1009,748)(-1009,742){3}
//: {4}(-1022,746)(-1022,658)(-1040,658){5}
wire G1;    //: /sn:0 {0}(-180,781)(-180,803)(-158,803)(-158,801){1}
wire w52;    //: /sn:0 {0}(-1324,-21)(-301,-21)(-301,397){1}
//: {2}(-299,399)(-279,399)(-279,381){3}
//: {4}(-301,401)(-301,443){5}
wire w17;    //: /sn:0 {0}(340,468)(340,444)(320,444)(320,405){1}
//: {2}(320,401)(320,345){3}
//: {4}(318,403)(306,403)(306,415)(291,415)(291,405){5}
wire w27;    //: /sn:0 {0}(-671,683)(-671,677)(-693,677)(-693,593){1}
//: {2}(-693,589)(-693,551){3}
//: {4}(-695,591)(-726,591)(-726,580){5}
wire w44;    //: /sn:0 {0}(-1368,841)(-1368,770){1}
//: {2}(-1368,766)(-1368,649)(-1387,649){3}
//: {4}(-1370,768)(-1388,768)(-1388,755){5}
wire w75;    //: /sn:0 {0}(-977,-377)(1505,-377)(1505,-36){1}
//: {2}(1507,-34)(1522,-34)(1522,-47){3}
//: {4}(1505,-32)(1505,-12)(1509,-12)(1509,1){5}
wire w35;    //: /sn:0 {0}(1028,243)(1028,172){1}
//: {2}(1028,168)(1028,51)(1009,51){3}
//: {4}(1026,170)(1008,170)(1008,157){5}
wire w33;    //: /sn:0 {0}(1305,243)(1305,210)(1374,210)(1374,152){1}
//: {2}(1376,150)(1387,150)(1387,144){3}
//: {4}(1374,148)(1374,60)(1356,60){5}
wire w28;    //: /sn:0 {0}(-1015,841)(-1015,808){1}
//: {2}(-1013,806)(-972,806)(-972,796){3}
//: {4}(-1015,804)(-1015,766)(-958,766)(-958,716){5}
wire w67;    //: /sn:0 {0}(-1225,-275)(190,-275)(190,184){1}
//: {2}(192,186)(199,186)(199,176){3}
//: {4}(190,188)(190,219){5}
wire w14;    //: /sn:0 {0}(-316,683)(-316,632){1}
//: {2}(-316,628)(-316,601)(-301,601)(-301,560){3}
//: {4}(-318,630)(-334,630)(-334,621){5}
wire w45;    //: /sn:0 {0}(-1214,658)(-1193,658)(-1193,779){1}
//: {2}(-1195,781)(-1207,781)(-1207,773){3}
//: {4}(-1193,783)(-1193,815)(-1226,815)(-1226,841){5}
wire S13;    //: /sn:0 {0}(-1429,749)(-1429,760)(-1415,760)(-1415,709){1}
wire w49;    //: /sn:0 {0}(-1431,25)(-967,25)(-967,577)(-948,577){1}
//: {2}(-946,575)(-946,572)(-929,572)(-929,555){3}
//: {4}(-946,579)(-946,599){5}
wire w69;    //: /sn:0 {0}(-1261,-261)(-81,-261)(-81,404){1}
//: {2}(-79,406)(-64,406)(-64,393){3}
//: {4}(-81,408)(-81,428)(-77,428)(-77,441){5}
wire P;    //: /sn:0 {0}(1333,341)(1333,370)(1361,370)(1361,360){1}
wire w11;    //: /sn:0 {0}(479,468)(479,417){1}
//: {2}(479,413)(479,386)(494,386)(494,345){3}
//: {4}(477,415)(461,415)(461,406){5}
wire w41;    //: /sn:0 {0}(-281,683)(-281,650)(-212,650)(-212,592){1}
//: {2}(-210,590)(-199,590)(-199,584){3}
//: {4}(-212,588)(-212,500)(-230,500){5}
wire w2;    //: /sn:0 {0}(-1503,56)(-1298,56)(-1298,550){1}
//: {2}(-1296,552)(-1281,552)(-1281,541){3}
//: {4}(-1298,554)(-1298,598)(-1297,598)(-1297,601){5}
wire w48;    //: /sn:0 {0}(-1467,42)(-1111,42)(-1111,555){1}
//: {2}(-1109,557)(-1089,557)(-1089,539){3}
//: {4}(-1111,559)(-1111,601){5}
wire w74;    //: /sn:0 {0}(-1083,-335)(981,-335)(981,-41){1}
//: {2}(983,-39)(990,-39)(990,-49){3}
//: {4}(981,-37)(981,-6){5}
wire w47;    //: /sn:0 {0}(-1536,881)(-1569,881)(-1569,821){1}
wire S12;    //: /sn:0 {0}(-877,716)(-877,782)(-859,782)(-859,774){1}
wire w15;    //: /sn:0 {0}(1131,243)(1131,219)(1111,219)(1111,180){1}
//: {2}(1111,176)(1111,120){3}
//: {4}(1109,178)(1097,178)(1097,190)(1082,190)(1082,180){5}
wire w5;    //: /sn:0 {0}(627,468)(627,462)(685,462)(685,427){1}
//: {2}(687,425)(695,425)(695,408){3}
//: {4}(685,423)(685,343){5}
wire w38;    //: /sn:0 {0}(514,468)(514,435)(583,435)(583,377){1}
//: {2}(585,375)(596,375)(596,369){3}
//: {4}(583,373)(583,285)(565,285){5}
wire P0;    //: /sn:0 {0}(542,566)(542,595)(570,595)(570,585){1}
wire w55;    //: /sn:0 {0}(-1218,-63)(307,-63)(307,177){1}
//: {2}(309,179)(324,179)(324,168){3}
//: {4}(307,181)(307,225)(308,225)(308,228){5}
wire w61;    //: /sn:0 {0}(-1005,-151)(1450,-151)(1450,-26){1}
//: {2}(1452,-24)(1467,-24)(1467,-43){3}
//: {4}(1450,-22)(1450,1){5}
wire S3;    //: /sn:0 {0}(967,151)(967,162)(981,162)(981,111){1}
wire w43;    //: /sn:0 {0}(-1481,841)(-1481,835)(-1503,835)(-1503,751){1}
//: {2}(-1503,747)(-1503,709){3}
//: {4}(-1505,749)(-1536,749)(-1536,738){5}
wire S14;    //: /sn:0 {0}(-1272,750)(-1272,757)(-1242,757)(-1242,718){1}
wire w64;    //: /sn:0 {0}(-1475,-170)(-1248,-170)(-1248,542){1}
//: {2}(-1246,544)(-1225,544)(-1225,533){3}
//: {4}(-1248,546)(-1248,583)(-1246,583)(-1246,601){5}
wire w9;    //: /sn:0 {0}(1270,243)(1270,192){1}
//: {2}(1270,188)(1270,161)(1285,161)(1285,120){3}
//: {4}(1268,190)(1252,190)(1252,181){5}
wire w26;    //: /sn:0 {0}(-618,683)(-618,677)(-648,677)(-648,620){1}
//: {2}(-648,616)(-648,551){3}
//: {4}(-650,618)(-669,618)(-669,607){5}
wire S10;    //: /sn:0 {0}(-462,592)(-462,599)(-432,599)(-432,560){1}
wire P2;    //: /sn:0 {0}(-1063,939)(-1063,968)(-1035,968)(-1035,958){1}
wire w76;    //: /sn:0 {0}(-1331,-231)(-438,-231)(-438,384){1}
//: {2}(-436,386)(-415,386)(-415,375){3}
//: {4}(-438,388)(-438,425)(-436,425)(-436,443){5}
wire S2;    //: /sn:0 {0}(1124,152)(1124,159)(1154,159)(1154,120){1}
wire w40;    //: /sn:0 {0}(-404,500)(-383,500)(-383,621){1}
//: {2}(-385,623)(-397,623)(-397,615){3}
//: {4}(-383,625)(-383,657)(-416,657)(-416,683){5}
wire S15;    //: /sn:0 {0}(-1087,746)(-1087,753)(-1068,753)(-1068,718){1}
wire w51;    //: /sn:0 {0}(-1359,-5)(-488,-5)(-488,392){1}
//: {2}(-486,394)(-471,394)(-471,383){3}
//: {4}(-488,396)(-488,440)(-487,440)(-487,443){5}
wire w57;    //: /sn:0 {0}(-1147,-94)(662,-94)(662,199){1}
//: {2}(664,201)(676,201)(676,182){3}
//: {4}(660,201)(659,201)(659,226){5}
wire w77;    //: /sn:0 {0}(-1190,-289)(357,-289)(357,169){1}
//: {2}(359,171)(380,171)(380,160){3}
//: {4}(357,173)(357,210)(359,210)(359,228){5}
//: enddecls

  CarryLookahead_Logic g4 (.G0(w3), .P0(w4), .G1(w9), .P1(w10), .G2(w15), .P2(w16), .G3(w21), .P3(w22), .Cin(w0), .C3(w35), .C2(w34), .C1(w33), .Cout(Cin0), .GG(G), .PG(P));   //: @(861, 244) /sz:(639, 96) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>0 Ti3>0 Ti4>0 Ti5>0 Ti6>0 Ti7>0 Ri0>9 To0<0 To1<5 To2<0 Lo0<7 Bo0<0 Bo1<0 ]
  //: joint g116 (w52) @(-301, 399) /w:[ 2 1 -1 4 ]
  //: switch g164 (w73) @(-1064,-349) /sn:0 /w:[ 0 ] /st:1
  //: switch g8 (w1) @(-1557,72) /sn:0 /w:[ 0 ] /st:0
  led g197 (.I(w29));   //: @(-1144,772) /sn:0 /w:[ 5 ] /type:0
  //: switch g157 (w68) @(-1171,-305) /sn:0 /w:[ 0 ] /st:1
  //: switch g17 (w48) @(-1484,42) /sn:0 /w:[ 0 ] /st:1
  led g258 (.I(w42));   //: @(-1479,758) /sn:0 /w:[ 5 ] /type:0
  led g224 (.I(w46));   //: @(-1009,735) /sn:0 /w:[ 3 ] /type:0
  CarryLookahead_Logic g137 (.G0(w7), .P0(w28), .G1(w29), .P1(w30), .G2(w31), .P2(w32), .G3(w42), .P3(w43), .Cin(Cin2), .C3(w44), .C2(w45), .C1(w46), .Cout(w47), .GG(G2), .PG(P2));   //: @(-1535, 842) /sz:(639, 96) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>0 Ti3>0 Ti4>0 Ti5>0 Ti6>0 Ti7>0 Ri0>0 To0<0 To1<5 To2<0 Lo0<0 Bo0<0 Bo1<0 ]
  //: joint g226 (w75) @(1505, -34) /w:[ 2 1 -1 4 ]
  //: switch g74 (w54) @(-1270,-49) /sn:0 /w:[ 0 ] /st:1
  led g92 (.I(w67));   //: @(199,169) /sn:0 /w:[ 3 ] /type:0
  led g30 (.I(w34));   //: @(1189,168) /sn:0 /w:[ 3 ] /type:0
  //: joint g198 (w46) @(-1022, 748) /w:[ 2 4 -1 1 ]
  //: switch g77 (w56) @(-1199,-79) /sn:0 /w:[ 0 ] /st:1
  //: joint g183 (w62) @(-891, 564) /w:[ 2 -1 1 4 ]
  //: joint g130 (w59) @(1098, -39) /w:[ -1 2 1 4 ]
  PFA_v1 g1 (.A(w70), .B(w60), .C(w33), .S(S1), .P(w10), .G(w9));   //: @(1229, 4) /sz:(126, 115) /sn:0 /p:[ Ti0>5 Ti1>5 Ri0>5 Bo0<1 Bo1<3 Bo2<3 ]
  led g214 (.I(w1));   //: @(-1453,556) /sn:0 /w:[ 3 ] /type:0
  //: joint g111 (w48) @(-1111, 557) /w:[ 2 1 -1 4 ]
  led g144 (.I(w68));   //: @(561,180) /sn:0 /w:[ 3 ] /type:0
  //: joint g51 (w22) @(893, 151) /w:[ -1 2 4 1 ]
  //: joint g179 (w64) @(-1248, 544) /w:[ 2 1 -1 4 ]
  led g260 (.I(w66));   //: @(-1044,553) /sn:0 /w:[ 3 ] /type:0
  led g190 (.I(w71));   //: @(-234,395) /sn:0 /w:[ 3 ] /type:0
  led g161 (.I(w25));   //: @(-540,617) /sn:0 /w:[ 5 ] /type:0
  //: joint g259 (w32) @(-1330, 798) /w:[ -1 2 4 1 ]
  led g70 (.I(w74));   //: @(990,-56) /sn:0 /w:[ 3 ] /type:0
  //: joint g206 (w43) @(-1503, 749) /w:[ -1 2 4 1 ]
  //: joint g103 (w17) @(320, 403) /w:[ -1 2 4 1 ]
  //: switch g65 (w53) @(-1306,-35) /sn:0 /w:[ 0 ] /st:0
  led g10 (.I(w14));   //: @(-334,614) /sn:0 /w:[ 5 ] /type:0
  led g25 (.I(S11));   //: @(-277,581) /sn:0 /w:[ 0 ] /type:0
  //: joint g149 (w20) @(-475, 618) /w:[ -1 2 4 1 ]
  //: joint g220 (w73) @(1148, -54) /w:[ 2 -1 1 4 ]
  led g64 (.I(w60));   //: @(1307,-66) /sn:0 /w:[ 3 ] /type:0
  led g185 (.I(S8));   //: @(-49,609) /sn:0 /w:[ 1 ] /type:0
  led g72 (.I(w58));   //: @(943,-42) /sn:0 /w:[ 3 ] /type:0
  //: joint g49 (w21) @(938, 178) /w:[ -1 2 4 1 ]
  led g251 (.I(S14));   //: @(-1272,743) /sn:0 /w:[ 0 ] /type:0
  led g142 (.I(w23));   //: @(126,385) /sn:0 /w:[ 5 ] /type:0
  //: joint g6 (w0) @(1596, 56) /w:[ 1 -1 2 4 ]
  //: joint g136 (w61) @(1450, -24) /w:[ 2 1 -1 4 ]
  led g7 (.I(Cin0));   //: @(827,216) /sn:0 /w:[ 9 ] /type:0
  led g56 (.I(w0));   //: @(1625,232) /sn:0 /w:[ 7 ] /type:0
  led g58 (.I(w75));   //: @(1522,-54) /sn:0 /w:[ 3 ] /type:0
  //: joint g124 (w56) @(494, 184) /w:[ 2 1 -1 4 ]
  //: joint g35 (w15) @(1111, 178) /w:[ -1 2 4 1 ]
  led g200 (.I(w45));   //: @(-1207,766) /sn:0 /w:[ 3 ] /type:0
  led g98 (.I(w54));   //: @(152,183) /sn:0 /w:[ 3 ] /type:0
  led g181 (.I(S10));   //: @(-462,585) /sn:0 /w:[ 0 ] /type:0
  //: joint g204 (w30) @(-1156, 763) /w:[ -1 2 4 1 ]
  //: joint g192 (w76) @(-438, 386) /w:[ 2 1 -1 4 ]
  led g85 (.I(S7));   //: @(518,366) /sn:0 /w:[ 0 ] /type:0
  led g67 (.I(w50));   //: @(-643,398) /sn:0 /w:[ 3 ] /type:0
  led g126 (.I(w17));   //: @(291,398) /sn:0 /w:[ 5 ] /type:0
  led g208 (.I(w63));   //: @(-1406,542) /sn:0 /w:[ 3 ] /type:0
  led g54 (.I(G));   //: @(1428,354) /sn:0 /w:[ 1 ] /type:0
  PFA_v1 g33 (.A(w71), .B(w52), .C(w41), .S(S11), .P(w19), .G(w14));   //: @(-357, 444) /sz:(126, 115) /sn:0 /p:[ Ti0>5 Ti1>5 Ri0>5 Bo0<1 Bo1<3 Bo2<3 ]
  led g40 (.I(S3));   //: @(967,144) /sn:0 /w:[ 0 ] /type:0
  led g52 (.I(P));   //: @(1361,353) /sn:0 /w:[ 1 ] /type:0
  led g81 (.I(w11));   //: @(461,399) /sn:0 /w:[ 5 ] /type:0
  //: joint g132 (w6) @(590, 433) /w:[ 2 4 -1 1 ]
  led g163 (.I(G1));   //: @(-158,794) /sn:0 /w:[ 1 ] /type:0
  led g108 (.I(w38));   //: @(596,362) /sn:0 /w:[ 3 ] /type:0
  //: joint g210 (w68) @(537, 197) /w:[ 2 1 -1 4 ]
  //: joint g12 (w41) @(-212, 590) /w:[ 2 4 -1 1 ]
  led g217 (.I(w47));   //: @(-1569,814) /sn:0 /w:[ 1 ] /type:0
  led g222 (.I(w2));   //: @(-1281,534) /sn:0 /w:[ 3 ] /type:0
  //: joint g131 (w5) @(685, 425) /w:[ 2 4 -1 1 ]
  led g106 (.I(w55));   //: @(324,161) /sn:0 /w:[ 3 ] /type:0
  //: joint g177 (w8) @(-110, 640) /w:[ 2 4 -1 1 ]
  PFA_v1 g194 (.A(w63), .B(w1), .C(w44), .S(S13), .P(w43), .G(w42));   //: @(-1514, 593) /sz:(126, 115) /sn:0 /p:[ Ti0>5 Ti1>5 Ri0>3 Bo0<1 Bo1<3 Bo2<3 ]
  led g96 (.I(w56));   //: @(516,159) /sn:0 /w:[ 3 ] /type:0
  //: joint g209 (w77) @(357, 171) /w:[ 2 1 -1 4 ]
  led g221 (.I(w62));   //: @(-874,544) /sn:0 /w:[ 3 ] /type:0
  led g117 (.I(G0));   //: @(637,579) /sn:0 /w:[ 1 ] /type:0
  //: joint g196 (w67) @(190, 186) /w:[ 2 1 -1 4 ]
  //: joint g114 (w51) @(-488, 394) /w:[ 2 1 -1 4 ]
  //: joint g19 (w3) @(1476, 200) /w:[ 2 4 -1 1 ]
  PFA_v1 g78 (.A(w67), .B(w54), .C(w36), .S(S5), .P(w24), .G(w23));   //: @(91, 220) /sz:(126, 115) /sn:0 /p:[ Ti0>5 Ti1>5 Ri0>3 Bo0<1 Bo1<3 Bo2<3 ]
  led g125 (.I(w12));   //: @(422,376) /sn:0 /w:[ 5 ] /type:0
  //: joint g219 (w31) @(-1285, 776) /w:[ -1 2 4 1 ]
  //: joint g155 (w40) @(-383, 623) /w:[ -1 1 2 4 ]
  led g105 (.I(w72));   //: @(731,171) /sn:0 /w:[ 3 ] /type:0
  //: joint g113 (w50) @(-661, 419) /w:[ -1 2 1 4 ]
  //: joint g223 (w70) @(1328, -28) /w:[ 2 1 -1 4 ]
  //: switch g93 (w59) @(-1092,-123) /sn:0 /w:[ 0 ] /st:0
  led g100 (.I(w24));   //: @(69,358) /sn:0 /w:[ 5 ] /type:0
  //: joint g63 (w26) @(-648, 618) /w:[ -1 2 4 1 ]
  led g212 (.I(w48));   //: @(-1089,532) /sn:0 /w:[ 3 ] /type:0
  led g205 (.I(w49));   //: @(-929,548) /sn:0 /w:[ 3 ] /type:0
  led g43 (.I(w53));   //: @(-119,390) /sn:0 /w:[ 3 ] /type:0
  led g38 (.I(w35));   //: @(1008,150) /sn:0 /w:[ 5 ] /type:0
  //: joint g211 (w72) @(714, 191) /w:[ 2 1 -1 4 ]
  //: joint g244 (Cin2) @(-759, 687) /w:[ -1 4 3 6 ]
  //: joint g215 (Cin2) @(-800, 664) /w:[ 2 8 -1 1 ]
  led g101 (.I(Cin1));   //: @(36,441) /sn:0 /w:[ 7 ] /type:0
  PFA_v1 g0 (.A(w75), .B(w61), .C(w0), .S(S0), .P(w4), .G(w3));   //: @(1420, 2) /sz:(126, 115) /sn:0 /p:[ Ti0>5 Ti1>5 Ri0>3 Bo0<0 Bo1<5 Bo2<5 ]
  led g48 (.I(w21));   //: @(917,160) /sn:0 /w:[ 5 ] /type:0
  //: joint g37 (w16) @(1066, 200) /w:[ -1 2 4 1 ]
  led g122 (.I(w77));   //: @(380,153) /sn:0 /w:[ 3 ] /type:0
  //: switch g80 (w58) @(-1128,-109) /sn:0 /w:[ 0 ] /st:0
  //: switch g95 (w61) @(-1022,-151) /sn:0 /w:[ 0 ] /st:1
  led g120 (.I(P0));   //: @(570,578) /sn:0 /w:[ 1 ] /type:0
  //: switch g76 (w55) @(-1235,-63) /sn:0 /w:[ 0 ] /st:0
  //: joint g189 (w25) @(-520, 640) /w:[ -1 2 4 1 ]
  //: joint g178 (w13) @(-205, 648) /w:[ 2 4 -1 1 ]
  //: switch g170 (w76) @(-1348,-231) /sn:0 /w:[ 0 ] /st:1
  //: switch g44 (w49) @(-1448,25) /sn:0 /w:[ 0 ] /st:0
  CarryLookahead_Logic g75 (.G0(w5), .P0(w6), .G1(w11), .P1(w12), .G2(w17), .P2(w18), .G3(w23), .P3(w24), .Cin(Cin0), .C3(w36), .C2(w37), .C1(w38), .Cout(Cin1), .GG(G0), .PG(P0));   //: @(70, 469) /sz:(639, 96) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>0 Ti3>0 Ti4>0 Ti5>0 Ti6>0 Ti7>0 Ri0>13 To0<0 To1<5 To2<0 Lo0<9 Bo0<0 Bo1<0 ]
  led g152 (.I(w51));   //: @(-471,376) /sn:0 /w:[ 3 ] /type:0
  //: joint g182 (w66) @(-1068, 570) /w:[ 2 1 -1 4 ]
  //: switch g159 (w70) @(-1029,-363) /sn:0 /w:[ 0 ] /st:1
  //: switch g47 (w50) @(-1411,10) /sn:0 /w:[ 0 ] /st:1
  //: switch g16 (w2) @(-1520,56) /sn:0 /w:[ 0 ] /st:0
  PFA_v1 g3 (.A(w74), .B(w58), .C(w35), .S(S3), .P(w22), .G(w21));   //: @(882, -5) /sz:(126, 115) /sn:0 /p:[ Ti0>5 Ti1>5 Ri0>3 Bo0<1 Bo1<3 Bo2<3 ]
  //: joint g90 (w24) @(102, 376) /w:[ -1 2 4 1 ]
  //: joint g109 (w37) @(412, 408) /w:[ -1 1 2 4 ]
  led g26 (.I(w9));   //: @(1252,174) /sn:0 /w:[ 5 ] /type:0
  //: joint g143 (w18) @(275, 425) /w:[ -1 2 4 1 ]
  //: joint g174 (Cin1) @(36, 498) /w:[ -1 6 5 8 ]
  //: joint g128 (Cin0) @(832, 283) /w:[ 6 -1 8 5 ]
  PFA_v1 g2 (.A(w73), .B(w59), .C(w34), .S(S2), .P(w16), .G(w15));   //: @(1055, 4) /sz:(126, 115) /sn:0 /p:[ Ti0>5 Ti1>5 Ri0>0 Bo0<1 Bo1<3 Bo2<3 ]
  //: switch g158 (w69) @(-1278,-261) /sn:0 /w:[ 0 ] /st:1
  led g91 (.I(w5));   //: @(695,401) /sn:0 /w:[ 3 ] /type:0
  //: joint g23 (w33) @(1374, 150) /w:[ 2 4 -1 1 ]
  //: joint g141 (w11) @(479, 415) /w:[ -1 2 4 1 ]
  //: joint g127 (Cin0) @(805, 477) /w:[ 1 2 -1 12 ]
  led g104 (.I(Cin0));   //: @(834,457) /sn:0 /w:[ 0 ] /type:0
  PFA_v1 g86 (.A(w68), .B(w56), .C(w38), .S(S7), .P(w12), .G(w11));   //: @(438, 229) /sz:(126, 115) /sn:0 /p:[ Ti0>5 Ti1>5 Ri0>5 Bo0<1 Bo1<3 Bo2<3 ]
  //: joint g39 (w35) @(1028, 170) /w:[ -1 2 4 1 ]
  led g24 (.I(S1));   //: @(1309,141) /sn:0 /w:[ 0 ] /type:0
  //: joint g29 (w10) @(1240, 165) /w:[ -1 2 4 1 ]
  //: joint g121 (w54) @(134, 201) /w:[ 2 1 -1 4 ]
  //: joint g110 (w2) @(-1298, 552) /w:[ 2 1 -1 4 ]
  led g60 (.I(w61));   //: @(1467,-50) /sn:0 /w:[ 3 ] /type:0
  led g250 (.I(w28));   //: @(-972,789) /sn:0 /w:[ 3 ] /type:0
  led g168 (.I(w76));   //: @(-415,368) /sn:0 /w:[ 3 ] /type:0
  PFA_v1 g199 (.A(w64), .B(w2), .C(w45), .S(S14), .P(w32), .G(w31));   //: @(-1341, 602) /sz:(126, 115) /sn:0 /p:[ Ti0>5 Ti1>5 Ri0>0 Bo0<1 Bo1<3 Bo2<3 ]
  led g18 (.I(w3));   //: @(1486,176) /sn:0 /w:[ 3 ] /type:0
  //: joint g257 (w29) @(-1126, 788) /w:[ -1 2 4 1 ]
  //: joint g82 (w38) @(583, 375) /w:[ 2 4 -1 1 ]
  //: joint g248 (w28) @(-1015, 806) /w:[ 2 4 -1 1 ]
  led g119 (.I(S5));   //: @(176,369) /sn:0 /w:[ 0 ] /type:0
  //: switch g94 (w60) @(-1057,-137) /sn:0 /w:[ 0 ] /st:1
  //: joint g173 (Cin1) @(10, 692) /w:[ 1 2 -1 12 ]
  led g154 (.I(w41));   //: @(-199,577) /sn:0 /w:[ 3 ] /type:0
  //: joint g107 (w1) @(-1471, 574) /w:[ 2 1 -1 4 ]
  led g166 (.I(P1));   //: @(-225,793) /sn:0 /w:[ 1 ] /type:0
  led g256 (.I(w44));   //: @(-1388,748) /sn:0 /w:[ 5 ] /type:0
  led g188 (.I(w26));   //: @(-669,600) /sn:0 /w:[ 5 ] /type:0
  PFA_v1 g184 (.A(w69), .B(w53), .C(Cin1), .S(S8), .P(w13), .G(w8));   //: @(-166, 442) /sz:(126, 115) /sn:0 /p:[ Ti0>5 Ti1>5 Ri0>11 Bo0<0 Bo1<5 Bo2<5 ]
  led g172 (.I(w20));   //: @(-504,613) /sn:0 /w:[ 5 ] /type:0
  led g216 (.I(w43));   //: @(-1536,731) /sn:0 /w:[ 5 ] /type:0
  led g50 (.I(w22));   //: @(860,133) /sn:0 /w:[ 5 ] /type:0
  //: joint g193 (w71) @(-258, 412) /w:[ 2 1 -1 4 ]
  led g73 (.I(Cin2));   //: @(-759,656) /sn:0 /w:[ 5 ] /type:0
  CarryLookahead_Logic g9 (.G0(w8), .P0(w13), .G1(w14), .P1(w19), .G2(w20), .P2(w25), .G3(w26), .P3(w27), .Cin(Cin1), .C3(w39), .C2(w40), .C1(w41), .Cout(Cin2), .GG(G1), .PG(P1));   //: @(-725, 684) /sz:(639, 96) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>0 Ti3>0 Ti4>0 Ti5>0 Ti6>0 Ti7>0 Ri0>13 To0<0 To1<5 To2<0 Lo0<7 Bo0<0 Bo1<0 ]
  //: joint g133 (w60) @(1285, -41) /w:[ 2 1 -1 4 ]
  led g68 (.I(w59));   //: @(1115,-64) /sn:0 /w:[ 3 ] /type:0
  led g186 (.I(w39));   //: @(-578,590) /sn:0 /w:[ 5 ] /type:0
  led g71 (.I(w27));   //: @(-726,573) /sn:0 /w:[ 5 ] /type:0
  //: switch g59 (w52) @(-1341,-21) /sn:0 /w:[ 0 ] /st:0
  //: joint g102 (w58) @(925, -24) /w:[ 2 1 -1 4 ]
  //: switch g169 (w75) @(-994,-377) /sn:0 /w:[ 0 ] /st:0
  //: joint g31 (w34) @(1203, 183) /w:[ -1 1 2 4 ]
  led g22 (.I(w33));   //: @(1387,137) /sn:0 /w:[ 3 ] /type:0
  //: joint g225 (w45) @(-1193, 781) /w:[ -1 1 2 4 ]
  //: joint g87 (w36) @(237, 395) /w:[ -1 2 4 1 ]
  led g231 (.I(w32));   //: @(-1350,775) /sn:0 /w:[ 5 ] /type:0
  led g180 (.I(w13));   //: @(-162,631) /sn:0 /w:[ 3 ] /type:0
  //: joint g99 (Cin0) @(805, 283) /w:[ 4 -1 10 3 ]
  PFA_v1 g83 (.A(w77), .B(w55), .C(w37), .S(S6), .P(w18), .G(w17));   //: @(264, 229) /sz:(126, 115) /sn:0 /p:[ Ti0>5 Ti1>5 Ri0>0 Bo0<1 Bo1<3 Bo2<3 ]
  //: joint g45 (w27) @(-693, 591) /w:[ -1 2 4 1 ]
  led g36 (.I(w16));   //: @(1046,177) /sn:0 /w:[ 5 ] /type:0
  //: joint g41 (w39) @(-558, 610) /w:[ -1 2 4 1 ]
  //: joint g203 (w44) @(-1368, 768) /w:[ -1 2 4 1 ]
  //: joint g69 (Cin1) @(10, 498) /w:[ 4 -1 10 3 ]
  //: switch g156 (w67) @(-1242,-275) /sn:0 /w:[ 0 ] /st:1
  PFA_v1 g138 (.A(w72), .B(w57), .C(Cin0), .S(S4), .P(w6), .G(w5));   //: @(629, 227) /sz:(126, 115) /sn:0 /p:[ Ti0>5 Ti1>5 Ri0>11 Bo0<0 Bo1<5 Bo2<5 ]
  //: joint g42 (w19) @(-346, 605) /w:[ -1 2 4 1 ]
  //: joint g213 (w42) @(-1458, 776) /w:[ -1 2 4 1 ]
  PFA_v1 g254 (.A(w62), .B(w49), .C(Cin2), .S(S12), .P(w28), .G(w7));   //: @(-976, 600) /sz:(126, 115) /sn:0 /p:[ Ti0>5 Ti1>5 Ri0>9 Bo0<0 Bo1<5 Bo2<5 ]
  //: switch g167 (w74) @(-1100,-335) /sn:0 /w:[ 0 ] /st:0
  led g66 (.I(w73));   //: @(1171,-72) /sn:0 /w:[ 3 ] /type:0
  led g151 (.I(w69));   //: @(-64,386) /sn:0 /w:[ 3 ] /type:0
  led g233 (.I(G2));   //: @(-968,952) /sn:0 /w:[ 1 ] /type:0
  //: joint g191 (w65) @(-605, 401) /w:[ 2 -1 1 4 ]
  //: switch g162 (w72) @(-1136,-320) /sn:0 /w:[ 0 ] /st:1
  //: switch g153 (w66) @(-1456,-184) /sn:0 /w:[ 0 ] /st:0
  //: switch g146 (w63) @(-1529,-154) /sn:0 /w:[ 0 ] /st:0
  led g242 (.I(w31));   //: @(-1314,771) /sn:0 /w:[ 5 ] /type:0
  led g28 (.I(w10));   //: @(1213,151) /sn:0 /w:[ 5 ] /type:0
  //: joint g57 (w0) @(1596, 252) /w:[ 6 5 -1 8 ]
  led g34 (.I(w15));   //: @(1082,173) /sn:0 /w:[ 5 ] /type:0
  led g46 (.I(w8));   //: @(-100,616) /sn:0 /w:[ 3 ] /type:0
  led g241 (.I(w30));   //: @(-1183,749) /sn:0 /w:[ 5 ] /type:0
  led g150 (.I(Cin1));   //: @(39,672) /sn:0 /w:[ 0 ] /type:0
  led g14 (.I(w40));   //: @(-397,608) /sn:0 /w:[ 3 ] /type:0
  PFA_v1 g11 (.A(w65), .B(w50), .C(w39), .S(S9), .P(w27), .G(w26));   //: @(-704, 435) /sz:(126, 115) /sn:0 /p:[ Ti0>5 Ti1>5 Ri0>3 Bo0<1 Bo1<3 Bo2<3 ]
  //: joint g118 (w53) @(-136, 416) /w:[ 2 1 -1 4 ]
  //: switch g5 (w0) @(1686,55) /sn:0 /R:2 /w:[ 0 ] /st:0
  led g84 (.I(w37));   //: @(398,393) /sn:0 /w:[ 3 ] /type:0
  //: joint g112 (w49) @(-946, 577) /w:[ -1 2 1 4 ]
  led g201 (.I(S15));   //: @(-1087,739) /sn:0 /w:[ 0 ] /type:0
  //: joint g187 (w14) @(-316, 630) /w:[ -1 2 4 1 ]
  //: joint g123 (w55) @(307, 179) /w:[ 2 1 -1 4 ]
  //: joint g21 (w4) @(1381, 208) /w:[ 2 4 -1 1 ]
  led g61 (.I(w52));   //: @(-279,374) /sn:0 /w:[ 3 ] /type:0
  led g255 (.I(S12));   //: @(-859,767) /sn:0 /w:[ 1 ] /type:0
  led g115 (.I(w18));   //: @(255,402) /sn:0 /w:[ 5 ] /type:0
  //: switch g79 (w57) @(-1164,-94) /sn:0 /w:[ 0 ] /st:0
  led g32 (.I(S2));   //: @(1124,145) /sn:0 /w:[ 0 ] /type:0
  led g20 (.I(w4));   //: @(1424,191) /sn:0 /w:[ 3 ] /type:0
  led g235 (.I(S13));   //: @(-1429,742) /sn:0 /w:[ 0 ] /type:0
  //: switch g145 (w62) @(-1420,-201) /sn:0 /w:[ 0 ] /st:1
  //: joint g176 (w63) @(-1415, 559) /w:[ 2 1 -1 4 ]
  //: switch g175 (w77) @(-1207,-289) /sn:0 /w:[ 0 ] /st:0
  //: joint g97 (w23) @(147, 403) /w:[ -1 2 4 1 ]
  led g134 (.I(w6));   //: @(633,416) /sn:0 /w:[ 3 ] /type:0
  led g236 (.I(P2));   //: @(-1035,951) /sn:0 /w:[ 1 ] /type:0
  //: joint g129 (w57) @(662, 201) /w:[ 2 1 4 -1 ]
  //: switch g148 (w65) @(-1383,-216) /sn:0 /w:[ 0 ] /st:0
  led g89 (.I(w57));   //: @(676,175) /sn:0 /w:[ 3 ] /type:0
  led g15 (.I(S0));   //: @(1537,169) /sn:0 /w:[ 1 ] /type:0
  PFA_v1 g202 (.A(w66), .B(w48), .C(w46), .S(S15), .P(w30), .G(w29));   //: @(-1167, 602) /sz:(126, 115) /sn:0 /p:[ Ti0>5 Ti1>5 Ri0>5 Bo0<1 Bo1<3 Bo2<3 ]
  //: joint g27 (w9) @(1270, 190) /w:[ -1 2 4 1 ]
  //: switch g147 (w64) @(-1492,-170) /sn:0 /w:[ 0 ] /st:0
  led g165 (.I(S9));   //: @(-619,584) /sn:0 /w:[ 0 ] /type:0
  //: joint g247 (w7) @(-920, 798) /w:[ 2 4 -1 1 ]
  led g171 (.I(w19));   //: @(-373,591) /sn:0 /w:[ 5 ] /type:0
  //: joint g218 (w74) @(981, -39) /w:[ 2 1 -1 4 ]
  //: switch g160 (w71) @(-1313,-247) /sn:0 /w:[ 0 ] /st:1
  led g62 (.I(w70));   //: @(1352,-45) /sn:0 /w:[ 3 ] /type:0
  led g238 (.I(w64));   //: @(-1225,526) /sn:0 /w:[ 3 ] /type:0
  //: joint g88 (w12) @(449, 390) /w:[ -1 2 4 1 ]
  //: joint g195 (w69) @(-81, 406) /w:[ 2 1 -1 4 ]
  //: switch g55 (w51) @(-1376,-5) /sn:0 /w:[ 0 ] /st:1
  led g207 (.I(w7));   //: @(-910,774) /sn:0 /w:[ 3 ] /type:0
  led g140 (.I(w36));   //: @(217,375) /sn:0 /w:[ 5 ] /type:0
  led g53 (.I(w65));   //: @(-596,384) /sn:0 /w:[ 3 ] /type:0
  PFA_v1 g13 (.A(w76), .B(w51), .C(w40), .S(S10), .P(w25), .G(w20));   //: @(-531, 444) /sz:(126, 115) /sn:0 /p:[ Ti0>5 Ti1>5 Ri0>0 Bo0<1 Bo1<3 Bo2<3 ]
  led g139 (.I(S4));   //: @(746,394) /sn:0 /w:[ 1 ] /type:0
  led g135 (.I(S6));   //: @(333,370) /sn:0 /w:[ 0 ] /type:0

endmodule
