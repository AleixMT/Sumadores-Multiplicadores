//: version "1.8.7"

module main;    //: root_module
wire w4;    //: /sn:0 {0}(213,201)(213,261)(241,261)(241,251){1}
wire w0;    //: /sn:0 {0}(194,-64)(248,-64)(248,10){1}
wire w1;    //: /sn:0 {0}(380,62)(390,62)(390,77)(342,77)(342,93)(332,93){1}
wire w2;    //: /sn:0 {0}(-9,55)(-9,97)(75,97){1}
wire w5;    //: /sn:0 {0}(82,-57)(143,-57)(143,10){1}
//: enddecls

  led g4 (.I(w2));   //: @(-9,48) /sn:0 /w:[ 0 ] /type:0
  //: switch g3 (w1) @(363,62) /sn:0 /w:[ 0 ] /st:1
  //: switch g2 (w0) @(177,-64) /sn:0 /w:[ 0 ] /st:1
  //: switch g1 (w5) @(65,-57) /sn:0 /w:[ 0 ] /st:1
  led g5 (.I(w4));   //: @(241,244) /sn:0 /w:[ 1 ] /type:0
  FA g0 (.B(w0), .A(w5), .Cin(w1), .Cout(w2), .S(w4));   //: @(76, 11) /sz:(255, 189) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<1 Bo0<0 ]

endmodule

module FA(S, Cout, Cin, B, A);
//: interface  /sz:(255, 189) /bd:[ Ti0>B(172/255) Ti1>A(67/255) Ri0>Cin(82/189) Lo0<Cout(86/189) Bo0<S(137/255) ]
input B;    //: /sn:0 {0}(171,166)(186,166)(186,140)(219,140){1}
//: {2}(223,140)(251,140){3}
//: {4}(221,142)(221,245)(392,245){5}
input A;    //: /sn:0 {0}(157,108)(185,108)(185,135)(198,135){1}
//: {2}(202,135)(251,135){3}
//: {4}(200,137)(200,240)(392,240){5}
input Cin;    //: /sn:0 {0}(182,222)(336,222)(336,188){1}
//: {2}(338,186)(348,186)(348,205)(379,205){3}
//: {4}(336,184)(336,161)(346,161){5}
output Cout;    //: /sn:0 /dp:1 {0}(477,235)(508,235)(508,213)(518,213){1}
output S;    //: /sn:0 /dp:1 {0}(367,159)(480,159)(480,152)(490,152){1}
wire w7;    //: /sn:0 {0}(413,243)(446,243)(446,237)(456,237){1}
wire w4;    //: /sn:0 {0}(400,208)(446,208)(446,232)(456,232){1}
wire w2;    //: /sn:0 {0}(272,138)(297,138){1}
//: {2}(301,138)(336,138)(336,156)(346,156){3}
//: {4}(299,140)(299,210)(379,210){5}
//: enddecls

  //: output g4 (S) @(487,152) /sn:0 /w:[ 1 ]
  and g8 (.I0(A), .I1(B), .Z(w7));   //: @(403,243) /sn:0 /delay:" 1" /w:[ 5 5 0 ]
  //: output g3 (Cout) @(515,213) /sn:0 /w:[ 1 ]
  //: input g2 (Cin) @(180,222) /sn:0 /w:[ 0 ]
  //: input g1 (B) @(169,166) /sn:0 /w:[ 0 ]
  //: joint g10 (w2) @(299, 138) /w:[ 2 -1 1 4 ]
  xor g6 (.I0(w2), .I1(Cin), .Z(S));   //: @(357,159) /sn:0 /delay:" 2" /w:[ 3 5 0 ]
  and g7 (.I0(Cin), .I1(w2), .Z(w4));   //: @(390,208) /sn:0 /delay:" 1" /w:[ 3 5 0 ]
  //: joint g9 (Cin) @(336, 186) /w:[ 2 4 -1 1 ]
  //: joint g12 (B) @(221, 140) /w:[ 2 -1 1 4 ]
  xor g5 (.I0(A), .I1(B), .Z(w2));   //: @(262,138) /sn:0 /delay:" 2" /w:[ 3 3 0 ]
  //: joint g11 (A) @(200, 135) /w:[ 2 -1 1 4 ]
  //: input g0 (A) @(155,108) /sn:0 /w:[ 0 ]
  or g13 (.I0(w4), .I1(w7), .Z(Cout));   //: @(467,235) /sn:0 /delay:" 1" /w:[ 1 1 0 ]

endmodule
