//: version "1.8.7"

module CarryLookahead_Logic(C2, P0, G0, P3, GG, G1, PG, P1, C3, C4, P2, C1, G3, Cin, G2);
//: interface  /sz:(639, 96) /bd:[ Ti0>G0(557/639) Ti1>P0(520/639) Ti2>G1(409/639) Ti3>P1(368/639) Ti4>G2(270/639) Ti5>P2(227/639) Ti6>G3(107/639) Ti7>P3(54/639) Ri0>Cin(46/96) To0<C3(167/639) To1<C2(309/639) To2<C1(444/639) Lo0<Cout(39/96) Bo0<GG(545/639) Bo1<PG(472/639) ]
input G2;    //: /sn:0 {0}(370,94)(370,89){1}
//: {2}(372,87)(391,87)(391,405){3}
//: {4}(393,407)(653,407){5}
//: {6}(391,409)(391,517){7}
//: {8}(393,519)(553,519){9}
//: {10}(391,521)(391,739)(567,739){11}
//: {12}(370,85)(370,76)(371,76)(371,69){13}
output GG;    //: /sn:0 /dp:1 {0}(692,765)(708,765)(708,763)(718,763){1}
input P1;    //: /sn:0 {0}(569,809)(259,809)(259,686){1}
//: {2}(261,684)(564,684){3}
//: {4}(257,684)(255,684)(255,627){5}
//: {6}(257,625)(560,625){7}
//: {8}(255,623)(255,584){9}
//: {10}(257,582)(555,582){11}
//: {12}(255,580)(255,447)(245,447){13}
//: {14}(243,445)(243,422){15}
//: {16}(245,420)(549,420){17}
//: {18}(243,418)(243,325)(233,325){19}
//: {20}(231,323)(231,293){21}
//: {22}(233,291)(537,291){23}
//: {24}(231,289)(231,73){25}
//: {26}(231,327)(231,330)(543,330){27}
//: {28}(243,449)(243,450)(552,450){29}
output C3;    //: /sn:0 /dp:1 {0}(674,409)(712,409)(712,405)(722,405){1}
output PG;    //: /sn:0 /dp:1 {0}(585,681)(671,681){1}
input G0;    //: /sn:0 {0}(569,814)(205,814)(205,589){1}
//: {2}(207,587)(555,587){3}
//: {4}(205,585)(205,422)(195,422){5}
//: {6}(193,420)(193,298){7}
//: {8}(195,296)(537,296){9}
//: {10}(193,294)(193,199){11}
//: {12}(195,197)(540,197){13}
//: {14}(193,195)(193,70){15}
//: {16}(193,424)(193,425)(549,425){17}
output C4;    //: /sn:0 /dp:1 {0}(686,553)(707,553)(707,545)(717,545){1}
output C2;    //: /sn:0 /dp:1 {0}(634,311)(642,311)(642,312)(652,312){1}
input Cin;    //: /sn:0 {0}(560,635)(83,635)(83,462){1}
//: {2}(85,460)(552,460){3}
//: {4}(83,458)(83,342){5}
//: {6}(85,340)(543,340){7}
//: {8}(83,338)(83,215){9}
//: {10}(85,213)(596,213){11}
//: {12}(83,211)(83,68){13}
input P3;    //: /sn:0 /dp:1 {0}(553,524)(433,524){1}
//: {2}(431,522)(431,64){3}
//: {4}(431,526)(431,542){5}
//: {6}(433,544)(556,544){7}
//: {8}(431,546)(431,570){9}
//: {10}(433,572)(555,572){11}
//: {12}(431,574)(431,613){13}
//: {14}(433,615)(560,615){15}
//: {16}(431,617)(431,672){17}
//: {18}(433,674)(564,674){19}
//: {20}(431,676)(431,732){21}
//: {22}(433,734)(567,734){23}
//: {24}(431,736)(431,765){25}
//: {26}(433,767)(569,767){27}
//: {28}(431,769)(431,799)(569,799){29}
input G1;    //: /sn:0 /dp:1 {0}(569,777)(279,777)(279,556){1}
//: {2}(281,554)(556,554){3}
//: {4}(279,552)(279,389){5}
//: {6}(281,387)(548,387){7}
//: {8}(279,385)(279,313){9}
//: {10}(281,311)(613,311){11}
//: {12}(279,309)(279,72){13}
input G3;    //: /sn:0 {0}(665,563)(492,563){1}
//: {2}(490,561)(490,63){3}
//: {4}(490,565)(490,763)(671,763){5}
output C1;    //: /sn:0 /dp:1 {0}(617,211)(626,211)(626,212)(636,212){1}
input P0;    //: /sn:0 {0}(564,689)(140,689)(140,632){1}
//: {2}(142,630)(560,630){3}
//: {4}(140,628)(140,457){5}
//: {6}(142,455)(552,455){7}
//: {8}(140,453)(140,337){9}
//: {10}(142,335)(543,335){11}
//: {12}(140,333)(140,204){13}
//: {14}(142,202)(540,202){15}
//: {16}(140,200)(140,69){17}
input P2;    //: /sn:0 /dp:1 {0}(548,382)(323,382){1}
//: {2}(321,380)(321,68){3}
//: {4}(321,384)(321,413){5}
//: {6}(323,415)(549,415){7}
//: {8}(321,417)(321,443){9}
//: {10}(323,445)(552,445){11}
//: {12}(321,447)(321,543){13}
//: {14}(319,545)(317,545)(317,575){15}
//: {16}(319,577)(555,577){17}
//: {18}(317,579)(317,618){19}
//: {20}(319,620)(560,620){21}
//: {22}(317,622)(317,674){23}
//: {24}(319,676)(329,676)(329,804)(569,804){25}
//: {26}(315,676)(305,676)(305,772)(569,772){27}
//: {28}(317,678)(317,679)(564,679){29}
//: {30}(321,547)(321,549)(556,549){31}
wire w6;    //: /sn:0 {0}(613,316)(574,316)(574,335)(564,335){1}
wire w4;    //: /sn:0 {0}(577,549)(620,549)(620,548)(665,548){1}
wire w3;    //: /sn:0 {0}(569,385)(643,385)(643,402)(653,402){1}
wire w0;    //: /sn:0 /dp:1 {0}(613,306)(568,306)(568,294)(558,294){1}
wire w12;    //: /sn:0 {0}(671,768)(600,768)(600,772)(590,772){1}
wire w1;    //: /sn:0 /dp:1 {0}(671,758)(598,758)(598,737)(588,737){1}
wire w8;    //: /sn:0 {0}(570,420)(643,420)(643,412)(653,412){1}
wire w17;    //: /sn:0 {0}(574,522)(655,522)(655,543)(665,543){1}
wire w14;    //: /sn:0 {0}(581,625)(642,625)(642,558)(665,558){1}
wire w11;    //: /sn:0 {0}(573,452)(650,452)(650,417)(653,417){1}
wire w15;    //: /sn:0 {0}(671,773)(618,773)(618,806)(590,806){1}
wire w5;    //: /sn:0 {0}(561,200)(586,200)(586,208)(596,208){1}
wire w9;    //: /sn:0 {0}(665,553)(633,553)(633,579)(576,579){1}
//: enddecls

  and g8 (.I0(P1), .I1(G0), .Z(w0));   //: @(548,294) /sn:0 /tech:unit /w:[ 23 9 1 ]
  or g4 (.I0(G0), .I1(P0), .Z(w5));   //: @(551,200) /sn:0 /tech:unit /w:[ 13 15 0 ]
  //: joint g44 (P1) @(243, 447) /w:[ 13 14 -1 28 ]
  or g16 (.I0(w0), .I1(G1), .I2(w6), .Z(C2));   //: @(624,311) /sn:0 /tech:unit /w:[ 0 11 0 0 ]
  and g3 (.I0(w5), .I1(Cin), .Z(C1));   //: @(607,211) /sn:0 /tech:unit /w:[ 1 11 0 ]
  //: joint g47 (P2) @(317, 577) /w:[ 16 15 -1 18 ]
  //: joint g26 (G0) @(193, 296) /w:[ 8 10 -1 7 ]
  //: output g17 (C2) @(649,312) /sn:0 /w:[ 1 ]
  //: input g2 (P0) @(140,67) /sn:0 /R:3 /w:[ 17 ]
  //: joint g30 (Cin) @(83, 340) /w:[ 6 8 -1 5 ]
  //: joint g23 (G1) @(279, 311) /w:[ 10 12 -1 9 ]
  //: joint g24 (P2) @(321, 382) /w:[ 1 2 -1 4 ]
  //: input g1 (G0) @(193,68) /sn:0 /R:3 /w:[ 15 ]
  //: joint g39 (P3) @(431, 524) /w:[ 1 2 -1 4 ]
  and g60 (.I0(P3), .I1(P2), .I2(G1), .Z(w12));   //: @(580,772) /sn:0 /w:[ 27 27 0 1 ]
  //: joint g29 (P0) @(140, 335) /w:[ 10 12 -1 9 ]
  or g51 (.I0(w17), .I1(w4), .I2(w9), .I3(w14), .I4(G3), .Z(C4));   //: @(676,553) /sn:0 /w:[ 1 1 0 1 0 0 ]
  or g70 (.I0(w1), .I1(G3), .I2(w12), .I3(w15), .Z(GG));   //: @(682,765) /sn:0 /w:[ 0 5 0 0 0 ]
  //: input g18 (P3) @(431,62) /sn:0 /R:3 /w:[ 3 ]
  //: joint g65 (P1) @(259, 684) /w:[ 2 -1 4 1 ]
  //: joint g25 (P1) @(231, 325) /w:[ 19 20 -1 26 ]
  and g10 (.I0(P1), .I1(P0), .I2(Cin), .Z(w6));   //: @(554,335) /sn:0 /tech:unit /w:[ 27 11 7 1 ]
  //: joint g64 (P3) @(431, 734) /w:[ 22 21 -1 24 ]
  //: output g72 (GG) @(715,763) /sn:0 /w:[ 1 ]
  //: joint g49 (P0) @(140, 455) /w:[ 6 8 -1 5 ]
  //: input g6 (G1) @(279,70) /sn:0 /R:3 /w:[ 13 ]
  //: joint g50 (Cin) @(83, 460) /w:[ 2 4 -1 1 ]
  //: joint g68 (P2) @(317, 676) /w:[ 24 23 26 28 ]
  //: output g58 (PG) @(668,681) /sn:0 /w:[ 1 ]
  //: joint g56 (P1) @(255, 625) /w:[ 6 8 -1 5 ]
  and g35 (.I0(P3), .I1(P2), .I2(P1), .I3(G0), .Z(w9));   //: @(566,579) /sn:0 /w:[ 11 17 11 3 1 ]
  //: joint g9 (G0) @(193, 197) /w:[ 12 14 -1 11 ]
  //: input g7 (P1) @(231,71) /sn:0 /R:3 /w:[ 25 ]
  //: joint g71 (G3) @(490, 563) /w:[ 1 2 -1 4 ]
  and g59 (.I0(P3), .I1(G2), .Z(w1));   //: @(578,737) /sn:0 /w:[ 23 11 1 ]
  or g31 (.I0(w3), .I1(G2), .I2(w8), .I3(w11), .Z(C3));   //: @(664,409) /sn:0 /w:[ 1 5 1 1 0 ]
  and g22 (.I0(P2), .I1(P1), .I2(P0), .I3(Cin), .Z(w11));   //: @(563,452) /sn:0 /w:[ 11 29 7 3 0 ]
  //: joint g67 (P3) @(431, 767) /w:[ 26 25 -1 28 ]
  //: joint g54 (P3) @(431, 615) /w:[ 14 13 -1 16 ]
  and g36 (.I0(P3), .I1(P2), .I2(P1), .I3(P0), .I4(Cin), .Z(w14));   //: @(571,625) /sn:0 /w:[ 15 21 7 3 0 0 ]
  //: output g33 (C3) @(719,405) /sn:0 /w:[ 1 ]
  //: joint g41 (G1) @(279, 387) /w:[ 6 8 -1 5 ]
  //: joint g45 (G0) @(193, 422) /w:[ 5 6 -1 16 ]
  //: joint g69 (G0) @(205, 587) /w:[ 2 4 -1 1 ]
  //: joint g40 (P2) @(321, 445) /w:[ 10 9 -1 12 ]
  //: joint g42 (P3) @(431, 544) /w:[ 6 5 -1 8 ]
  //: output g52 (C4) @(714,545) /sn:0 /w:[ 1 ]
  //: joint g66 (G1) @(279, 554) /w:[ 2 4 -1 1 ]
  //: input g12 (P2) @(321,66) /sn:0 /R:3 /w:[ 3 ]
  //: joint g57 (P0) @(140, 630) /w:[ 2 4 -1 1 ]
  and g34 (.I0(P3), .I1(P2), .I2(G1), .Z(w4));   //: @(567,549) /sn:0 /w:[ 7 31 3 0 ]
  //: joint g28 (P1) @(243, 420) /w:[ 16 18 -1 15 ]
  //: joint g46 (P3) @(431, 572) /w:[ 10 9 -1 12 ]
  //: joint g14 (P0) @(140, 202) /w:[ 14 16 -1 13 ]
  //: joint g11 (Cin) @(83, 213) /w:[ 10 12 -1 9 ]
  //: output g5 (C1) @(633,212) /sn:0 /w:[ 1 ]
  and g61 (.I0(P3), .I1(P2), .I2(P1), .I3(G0), .Z(w15));   //: @(580,806) /sn:0 /w:[ 29 25 0 0 1 ]
  and g21 (.I0(P2), .I1(P1), .I2(G0), .Z(w8));   //: @(560,420) /sn:0 /w:[ 7 17 17 0 ]
  //: input g19 (G3) @(490,61) /sn:0 /R:3 /w:[ 3 ]
  //: joint g32 (G2) @(370, 87) /w:[ 2 12 -1 1 ]
  and g20 (.I0(P2), .I1(G1), .Z(w3));   //: @(559,385) /sn:0 /w:[ 0 7 0 ]
  //: joint g63 (G2) @(391, 519) /w:[ 8 7 -1 10 ]
  //: joint g38 (G2) @(391, 407) /w:[ 4 3 -1 6 ]
  //: joint g15 (P1) @(231, 291) /w:[ 22 24 -1 21 ]
  //: input g0 (Cin) @(83,66) /sn:0 /R:3 /w:[ 13 ]
  //: joint g43 (P2) @(321, 545) /w:[ -1 13 14 30 ]
  //: joint g27 (P2) @(321, 415) /w:[ 6 5 -1 8 ]
  //: joint g48 (P1) @(255, 582) /w:[ 10 12 -1 9 ]
  //: joint g62 (P3) @(431, 674) /w:[ 18 17 -1 20 ]
  and g37 (.I0(G2), .I1(P3), .Z(w17));   //: @(564,522) /sn:0 /w:[ 9 0 0 ]
  //: joint g55 (P2) @(317, 620) /w:[ 20 19 -1 22 ]
  and g53 (.I0(P3), .I1(P2), .I2(P1), .I3(P0), .Z(PG));   //: @(575,681) /sn:0 /w:[ 19 29 3 0 0 ]
  //: input g13 (G2) @(371,67) /sn:0 /R:3 /w:[ 13 ]

endmodule

module CLA_Adder_4bit(P, G);
//: interface  /sz:(209, 138) /bd:[ Ti0>A0(190/209) Ti1>A1(172/209) Ti2>A2(151/209) Ti3>A3(130/209) Ti4>B0(99/209) Ti5>B1(79/209) Ti6>B2(63/209) Ti7>B3(42/209) Ri0>Cin(59/138) Bo0<P(192/209) Bo1<G(148/209) ]
output G;    //: /sn:0 {0}(887,612)(887,656){1}
output P;    //: /sn:0 {0}(814,612)(814,660){1}
wire w16;    //: /sn:0 {0}(547,391)(547,457){1}
//: {2}(549,459)(579,459)(579,457){3}
//: {4}(547,461)(547,506)(569,506)(569,514){5}
wire w34;    //: /sn:0 {0}(651,514)(651,486)(684,486)(684,331)(677,331){1}
//: {2}(675,329)(675,319)(674,319)(674,308){3}
//: {4}(673,331)(663,331){5}
wire w25;    //: /sn:0 {0}(915,255)(925,255)(925,272){1}
wire w4;    //: /sn:0 {0}(922,389)(922,441)(863,441)(863,460){1}
//: {2}(865,462)(888,462)(888,474)(903,474)(903,464){3}
//: {4}(863,464)(863,501)(862,501)(862,514){5}
wire w0;    //: /sn:0 {0}(790,424)(790,434)(809,434)(809,391){1}
wire w22;    //: /sn:0 {0}(374,382)(374,428){1}
//: {2}(376,430)(400,430)(400,423){3}
//: {4}(374,432)(374,506)(396,506)(396,514){5}
wire w3;    //: /sn:0 {0}(960,389)(960,422)(958,422)(958,455){1}
//: {2}(960,457)(1026,457)(1026,491)(1042,491)(1042,481){3}
//: {4}(958,459)(958,506)(899,506)(899,514){5}
wire w20;    //: /sn:0 {0}(728,247)(731,247)(731,274){1}
wire w19;    //: /sn:0 {0}(608,253)(618,253)(618,274){1}
wire w18;    //: /sn:0 {0}(552,248)(557,248)(557,274){1}
wire w23;    //: /sn:0 {0}(462,382)(462,430)(478,430)(478,420){1}
wire w10;    //: /sn:0 {0}(721,391)(721,439){1}
//: {2}(723,441)(739,441)(739,428){3}
//: {4}(721,443)(721,474)(710,474)(710,514){5}
wire w24;    //: /sn:0 {0}(779,241)(792,241)(792,274){1}
wire w21;    //: /sn:0 {0}(419,382)(419,461){1}
//: {2}(421,463)(455,463)(455,449){3}
//: {4}(419,465)(419,506)(449,506)(449,514){5}
wire w1;    //: /sn:0 {0}(990,430)(990,440)(1003,440)(1003,389){1}
wire w32;    //: /sn:0 {0}(982,561)(1077,561)(1077,329){1}
//: {2}(1077,325)(1077,298)(1066,298){3}
//: {4}(1075,327)(1039,327)(1039,329)(1031,329){5}
wire w8;    //: /sn:0 {0}(369,234)(384,234)(384,265){1}
wire w17;    //: /sn:0 {0}(635,391)(635,435)(655,435)(655,425){1}
wire w33;    //: /sn:0 {0}(786,514)(786,479)(855,479)(855,333){1}
//: {2}(855,329)(855,319)(849,319)(849,289){3}
//: {4}(853,331)(837,331){5}
wire w35;    //: /sn:0 {0}(509,514)(509,335)(507,335)(507,324){1}
//: {2}(507,320)(507,310)(501,310)(501,277){3}
//: {4}(505,322)(490,322){5}
wire w14;    //: /sn:0 {0}(436,234)(445,234)(445,265){1}
wire w2;    //: /sn:0 {0}(309,520)(309,554)(341,554){1}
wire w15;    //: /sn:0 {0}(592,391)(592,432){1}
//: {2}(594,434)(608,434)(608,441)(623,441)(623,431){3}
//: {4}(592,436)(592,488)(612,488)(612,514){5}
wire w26;    //: /sn:0 {0}(972,248)(986,248)(986,272){1}
wire w9;    //: /sn:0 {0}(766,391)(766,434)(752,434)(752,469){1}
//: {2}(754,471)(760,471)(760,484)(775,484)(775,474){3}
//: {4}(752,473)(752,505)(751,505)(751,514){5}
//: enddecls

  CarryLookahead_Logic g4 (.G0(w3), .P0(w4), .G1(w9), .P1(w10), .G2(w15), .P2(w16), .G3(w21), .P3(w22), .Cin(w32), .C3(w35), .C2(w34), .C1(w33), .Cout(w2), .GG(G), .PG(P));   //: @(342, 515) /sz:(639, 96) /sn:0 /p:[ Ti0>5 Ti1>5 Ti2>5 Ti3>5 Ti4>5 Ti5>5 Ti6>5 Ti7>5 Ri0>0 To0<0 To1<0 To2<0 Lo0<1 Bo0<0 Bo1<0 ]
  //: switch g8 (w8) @(352,234) /sn:0 /w:[ 0 ] /st:1
  PFA_v1 g3 (.A(w8), .B(w14), .C(w35), .S(w23), .P(w22), .G(w21));   //: @(363, 266) /sz:(126, 115) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>5 Bo0<0 Bo1<0 Bo2<0 ]
  led g16 (.I(w33));   //: @(849,282) /sn:0 /w:[ 3 ] /type:0
  led g26 (.I(w3));   //: @(1042,474) /sn:0 /w:[ 3 ] /type:0
  //: joint g17 (w33) @(855, 331) /w:[ -1 2 4 1 ]
  PFA_v1 g2 (.A(w18), .B(w19), .C(w34), .S(w17), .P(w16), .G(w15));   //: @(536, 275) /sz:(126, 115) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>5 Bo0<0 Bo1<0 Bo2<0 ]
  led g30 (.I(w9));   //: @(775,467) /sn:0 /w:[ 3 ] /type:0
  led g23 (.I(w17));   //: @(655,418) /sn:0 /w:[ 1 ] /type:0
  //: joint g39 (w21) @(419, 463) /w:[ 2 1 -1 4 ]
  PFA_v1 g1 (.A(w20), .B(w24), .C(w33), .S(w0), .P(w10), .G(w9));   //: @(710, 275) /sz:(126, 115) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>5 Bo0<1 Bo1<0 Bo2<0 ]
  led g24 (.I(w0));   //: @(790,417) /sn:0 /w:[ 0 ] /type:0
  //: joint g29 (w4) @(863, 462) /w:[ 2 1 -1 4 ]
  led g18 (.I(w34));   //: @(674,301) /sn:0 /w:[ 3 ] /type:0
  //: switch g10 (w18) @(535,248) /sn:0 /w:[ 0 ] /st:1
  led g25 (.I(w1));   //: @(990,423) /sn:0 /w:[ 0 ] /type:0
  //: joint g6 (w32) @(1077, 327) /w:[ -1 2 4 1 ]
  //: joint g35 (w15) @(592, 434) /w:[ 2 1 -1 4 ]
  led g7 (.I(w2));   //: @(309,513) /sn:0 /w:[ 0 ] /type:0
  //: switch g9 (w14) @(419,234) /sn:0 /w:[ 0 ] /st:1
  //: joint g31 (w9) @(752, 471) /w:[ 2 1 -1 4 ]
  led g22 (.I(w23));   //: @(478,413) /sn:0 /w:[ 1 ] /type:0
  //: joint g41 (w22) @(374, 430) /w:[ 2 1 -1 4 ]
  led g36 (.I(w16));   //: @(579,450) /sn:0 /w:[ 3 ] /type:0
  //: joint g33 (w10) @(721, 441) /w:[ 2 1 -1 4 ]
  led g40 (.I(w22));   //: @(400,416) /sn:0 /w:[ 3 ] /type:0
  //: output g42 (P) @(814,657) /sn:0 /R:3 /w:[ 1 ]
  //: switch g12 (w20) @(711,247) /sn:0 /w:[ 0 ] /st:0
  led g34 (.I(w15));   //: @(623,424) /sn:0 /w:[ 3 ] /type:0
  led g28 (.I(w4));   //: @(903,457) /sn:0 /w:[ 3 ] /type:0
  //: switch g5 (w32) @(1049,298) /sn:0 /w:[ 3 ] /st:1
  //: switch g11 (w19) @(591,253) /sn:0 /w:[ 0 ] /st:0
  //: switch g14 (w25) @(898,255) /sn:0 /w:[ 0 ] /st:0
  //: joint g19 (w34) @(675, 331) /w:[ 1 2 4 -1 ]
  //: joint g21 (w35) @(507, 322) /w:[ -1 2 4 1 ]
  led g32 (.I(w10));   //: @(739,421) /sn:0 /w:[ 3 ] /type:0
  led g20 (.I(w35));   //: @(501,270) /sn:0 /w:[ 3 ] /type:0
  led g38 (.I(w21));   //: @(455,442) /sn:0 /w:[ 3 ] /type:0
  PFA_v1 g0 (.A(w25), .B(w26), .C(w32), .S(w1), .P(w4), .G(w3));   //: @(904, 273) /sz:(126, 115) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>5 Bo0<1 Bo1<0 Bo2<0 ]
  //: switch g15 (w26) @(955,248) /sn:0 /w:[ 0 ] /st:1
  //: output g43 (G) @(887,653) /sn:0 /R:3 /w:[ 1 ]
  //: joint g27 (w3) @(958, 457) /w:[ 2 1 -1 4 ]
  //: joint g37 (w16) @(547, 459) /w:[ 2 1 -1 4 ]
  //: switch g13 (w24) @(762,241) /sn:0 /w:[ 0 ] /st:1

endmodule

module PFA_v1(C, B, P, S, A, G);
//: interface  /sz:(126, 115) /bd:[ Ti0>A(21/126) Ti1>B(82/126) Ri0>C(56/115) Bo0<S(99/126) Bo1<P(11/126) Bo2<G(56/126) ]
input B;    //: /sn:0 {0}(144,200)(161,200){1}
//: {2}(165,200)(202,200)(202,177)(210,177){3}
//: {4}(163,202)(163,320){5}
//: {6}(165,322)(231,322){7}
//: {8}(163,324)(163,361)(240,361){9}
input A;    //: /sn:0 {0}(151,147)(178,147){1}
//: {2}(182,147)(202,147)(202,172)(210,172){3}
//: {4}(180,149)(180,317)(188,317){5}
//: {6}(192,317)(231,317){7}
//: {8}(190,319)(190,356)(240,356){9}
output G;    //: /sn:0 /dp:1 {0}(261,359)(337,359)(337,385)(346,385){1}
input C;    //: /sn:0 {0}(149,271)(266,271)(266,186)(276,186){1}
output P;    //: /sn:0 /dp:1 {0}(252,320)(312,320)(312,319)(322,319){1}
output S;    //: /sn:0 /dp:1 {0}(297,184)(394,184)(394,198)(406,198){1}
wire w2;    //: /sn:0 {0}(231,175)(267,175)(267,181)(276,181){1}
//: enddecls

  xor g4 (.I0(w2), .I1(C), .Z(S));   //: @(287,184) /sn:0 /delay:" 2" /w:[ 1 1 0 ]
  //: joint g8 (B) @(163, 200) /w:[ 2 -1 1 4 ]
  xor g3 (.I0(A), .I1(B), .Z(w2));   //: @(221,175) /sn:0 /delay:" 2" /w:[ 3 3 0 ]
  //: input g2 (C) @(147,271) /sn:0 /w:[ 0 ]
  //: input g1 (B) @(142,200) /sn:0 /w:[ 0 ]
  and g10 (.I0(A), .I1(B), .Z(G));   //: @(251,359) /sn:0 /delay:" 1" /w:[ 9 9 0 ]
  or g6 (.I0(A), .I1(B), .Z(P));   //: @(242,320) /sn:0 /delay:" 1" /w:[ 7 7 0 ]
  //: joint g7 (A) @(180, 147) /w:[ 2 -1 1 4 ]
  //: output g9 (P) @(319,319) /sn:0 /w:[ 1 ]
  //: joint g12 (A) @(190, 317) /w:[ 6 -1 5 8 ]
  //: output g5 (S) @(403,198) /sn:0 /w:[ 1 ]
  //: joint g11 (B) @(163, 322) /w:[ 6 5 -1 8 ]
  //: input g0 (A) @(149,147) /sn:0 /w:[ 0 ]
  //: output g13 (G) @(343,385) /sn:0 /w:[ 1 ]

endmodule

module main;    //: root_module
wire w13;    //: /sn:0 {0}(254,353)(254,363){1}
wire w6;    //: /sn:0 {0}(347,353)(347,363){1}
wire w16;    //: /sn:0 {0}(5,507)(5,587)(-85,587)(-85,681){1}
wire w7;    //: /sn:0 {0}(326,353)(326,363){1}
wire w58;    //: /sn:0 {0}(92,779)(92,807)(101,807)(101,817){1}
wire w34;    //: /sn:0 {0}(-636,374)(-636,364){1}
wire w4;    //: /sn:0 {0}(12,367)(12,357){1}
wire w39;    //: /sn:0 {0}(-527,374)(-527,364){1}
wire w56;    //: /sn:0 {0}(-464,721)(-454,721){1}
wire w0;    //: /sn:0 {0}(-76,367)(-76,357){1}
wire w3;    //: /sn:0 {0}(-19,367)(-19,357){1}
wire w22;    //: /sn:0 {0}(-256,374)(-256,364){1}
wire w36;    //: /sn:0 {0}(-600,374)(-600,364){1}
wire w20;    //: /sn:0 {0}(-308,374)(-308,364){1}
wire w30;    //: /sn:0 {0}(294,503)(294,632)(67,632)(67,681){1}
wire w37;    //: /sn:0 {0}(-569,374)(-569,364){1}
wire w42;    //: /sn:0 {0}(-551,514)(-551,643)(-346,643)(-346,681){1}
wire w12;    //: /sn:0 {0}(274,353)(274,363){1}
wire w18;    //: /sn:0 {0}(-344,374)(-344,364){1}
wire w19;    //: /sn:0 {0}(-328,374)(-328,364){1}
wire w10;    //: /sn:0 {0}(72,367)(72,357){1}
wire w23;    //: /sn:0 {0}(-235,374)(-235,364){1}
wire w54;    //: /sn:0 {0}(-144,681)(-144,434)(-197,434){1}
wire w21;    //: /sn:0 {0}(-277,374)(-277,364){1}
wire w24;    //: /sn:0 {0}(-217,374)(-217,364){1}
wire w31;    //: /sn:0 {0}(323,503)(323,655)(104,655)(104,681){1}
wire w1;    //: /sn:0 {0}(-55,367)(-55,357){1}
wire w32;    //: /sn:0 {0}(-289,514)(-289,630)(-226,630)(-226,681){1}
wire w53;    //: /sn:0 {0}(-9,681)(-9,654)(48,654)(48,561)(159,561)(159,427)(92,427){1}
wire w8;    //: /sn:0 {0}(33,367)(33,357){1}
wire w52;    //: /sn:0 {0}(187,728)(456,728)(456,425){1}
//: {2}(458,423)(489,423)(489,433)(497,433){3}
//: {4}(454,423)(385,423){5}
wire w27;    //: /sn:0 {0}(238,353)(238,363){1}
wire w17;    //: /sn:0 {0}(-365,374)(-365,364){1}
wire w28;    //: /sn:0 {0}(217,353)(217,363){1}
wire w33;    //: /sn:0 {0}(-657,374)(-657,364){1}
wire w35;    //: /sn:0 {0}(-620,374)(-620,364){1}
wire w11;    //: /sn:0 {0}(305,353)(305,363){1}
wire w2;    //: /sn:0 {0}(-39,367)(-39,357){1}
wire w15;    //: /sn:0 {0}(30,507)(30,619)(-44,619)(-44,681){1}
wire w5;    //: /sn:0 {0}(365,353)(365,363){1}
wire w38;    //: /sn:0 {0}(-548,374)(-548,364){1}
wire w55;    //: /sn:0 {0}(-309,681)(-309,616)(-450,616)(-450,434)(-489,434){1}
wire w43;    //: /sn:0 {0}(-583,514)(-583,671)(-399,671)(-399,681){1}
wire w9;    //: /sn:0 {0}(54,367)(54,357){1}
wire w26;    //: /sn:0 {0}(-259,514)(-259,603)(-183,603)(-183,681){1}
wire w40;    //: /sn:0 {0}(-509,374)(-509,364){1}
wire w57;    //: /sn:0 {0}(19,779)(19,810)(21,810)(21,820){1}
//: enddecls

  led g4 (.I(w58));   //: @(101,824) /sn:0 /R:2 /w:[ 1 ] /type:0
  CarryLookahead_Logic g3 (.G0(w31), .P0(w30), .G1(w15), .P1(w16), .G2(w26), .P2(w32), .G3(w42), .P3(w43), .Cin(w52), .C3(w55), .C2(w54), .C1(w53), .Cout(w56), .GG(w58), .PG(w57));   //: @(-453, 682) /sz:(639, 96) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Ti3>1 Ti4>1 Ti5>1 Ti6>1 Ti7>1 Ri0>0 To0<0 To1<0 To2<0 Lo0<1 Bo0<0 Bo1<0 ]
  CLA_Adder_4bit g2 (.A0(w40), .A1(w39), .A2(w38), .A3(w37), .B0(w36), .B1(w35), .B2(w34), .B3(w33), .Cin(w55), .P(w43), .G(w42));   //: @(-699, 375) /sz:(209, 138) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>0 Ti3>0 Ti4>0 Ti5>0 Ti6>0 Ti7>0 Ri0>1 Bo0<0 Bo1<0 ]
  CLA_Adder_4bit g1 (.A0(w24), .A1(w23), .A2(w22), .A3(w21), .B0(w20), .B1(w19), .B2(w18), .B3(w17), .Cin(w54), .P(w32), .G(w26));   //: @(-407, 375) /sz:(209, 138) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>0 Ti3>0 Ti4>0 Ti5>0 Ti6>0 Ti7>0 Ri0>1 Bo0<0 Bo1<0 ]
  //: switch g6 (w52) @(515,433) /sn:0 /R:2 /w:[ 3 ] /st:0
  //: joint g7 (w52) @(456, 423) /w:[ 2 -1 4 1 ]
  CLA_Adder_4bit g42 (.B3(w28), .B2(w27), .B1(w13), .B0(w12), .A3(w11), .A2(w7), .A1(w6), .A0(w5), .Cin(w52), .G(w31), .P(w30));   //: @(175, 364) /sz:(209, 138) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Ti3>1 Ti4>1 Ti5>1 Ti6>1 Ti7>1 Ri0>5 Bo0<0 Bo1<0 ]
  led g5 (.I(w57));   //: @(21,827) /sn:0 /R:2 /w:[ 1 ] /type:0
  CLA_Adder_4bit g0 (.A0(w10), .A1(w9), .A2(w8), .A3(w4), .B0(w3), .B1(w2), .B2(w1), .B3(w0), .Cin(w53), .P(w16), .G(w15));   //: @(-118, 368) /sz:(209, 138) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>0 Ti3>0 Ti4>0 Ti5>0 Ti6>0 Ti7>0 Ri0>1 Bo0<0 Bo1<0 ]

endmodule
