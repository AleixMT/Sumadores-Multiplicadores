//: version "1.8.7"

module CPA(C0, A1, S0, B2, A2, B3, S2, S3, A0, C4, B0, B1, A3, S1);
//: interface  /sz:(223, 91) /bd:[ Ti0>A3(11/223) Ti1>B3(29/223) Ti2>A2(48/223) Ti3>B2(66/223) Ti4>A1(83/223) Ti5>B1(103/223) Ti6>A0(118/223) Ti7>B0(136/223) Ri0>C0(34/91) Lo0<C4(39/91) Bo0<S0(175/223) Bo1<S1(127/223) Bo2<S2(76/223) Bo3<S3(39/223) ]
input A0;    //: /sn:0 {0}(709,242)(709,291)(707,291)(707,322){1}
output S1;    //: /sn:0 /dp:1 {0}(607,430)(607,503)(605,503)(605,506){1}
input C0;    //: /sn:0 {0}(847,365)(801,365){1}
input A3;    //: /sn:0 {0}(308,253)(308,290)(310,290)(310,331){1}
input A2;    //: /sn:0 {0}(448,236)(448,324)(447,324)(447,325){1}
input B2;    //: /sn:0 {0}(491,237)(491,325){1}
output C4;    //: /sn:0 {0}(217,374)(284,374){1}
input B1;    //: /sn:0 {0}(622,241)(622,310)(621,310)(621,320){1}
output S0;    //: /sn:0 /dp:1 {0}(748,422)(748,440)(749,440)(749,511){1}
input A1;    //: /sn:0 {0}(578,242)(578,320){1}
input B3;    //: /sn:0 {0}(352,249)(352,326)(351,326)(351,331){1}
output S3;    //: /sn:0 {0}(326,497)(326,456)(337,456)(337,426){1}
input B0;    //: /sn:0 {0}(761,241)(761,312)(763,312)(763,322){1}
output S2;    //: /sn:0 /dp:1 {0}(476,429)(476,497){1}
wire w6;    //: /sn:0 {0}(657,367)(688,367){1}
wire w4;    //: /sn:0 {0}(527,370)(550,370){1}
wire w3;    //: /sn:0 {0}(384,372)(419,372){1}
//: enddecls

  //: input g8 (C0) @(849,365) /sn:0 /R:2 /w:[ 0 ]
  //: input g4 (A1) @(578,240) /sn:0 /R:3 /w:[ 0 ]
  //: output g13 (S0) @(749,508) /sn:0 /R:3 /w:[ 1 ]
  //: input g3 (B2) @(491,235) /sn:0 /R:3 /w:[ 0 ]
  //: input g2 (A2) @(448,234) /sn:0 /R:3 /w:[ 0 ]
  //: input g1 (B3) @(352,247) /sn:0 /R:3 /w:[ 0 ]
  //: output g11 (S2) @(476,494) /sn:0 /R:3 /w:[ 1 ]
  FA g16 (.A(A1), .B(B1), .Cin(w6), .Cout(w4), .S(S1));   //: @(551, 321) /sz:(105, 108) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  //: output g10 (S3) @(326,494) /sn:0 /R:3 /w:[ 0 ]
  //: input g6 (A0) @(709,240) /sn:0 /R:3 /w:[ 0 ]
  //: output g9 (C4) @(220,374) /sn:0 /R:2 /w:[ 0 ]
  //: input g7 (B0) @(761,239) /sn:0 /R:3 /w:[ 0 ]
  FA g15 (.A(A2), .B(B2), .Cin(w4), .Cout(w3), .S(S2));   //: @(420, 326) /sz:(106, 102) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  FA g17 (.A(A0), .B(B0), .Cin(C0), .Cout(w6), .S(S0));   //: @(689, 323) /sz:(111, 98) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<1 Bo0<0 ]
  //: input g5 (B1) @(622,239) /sn:0 /R:3 /w:[ 0 ]
  FA g14 (.A(A3), .B(B3), .Cin(w3), .Cout(C4), .S(S3));   //: @(285, 332) /sz:(98, 93) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<1 ]
  //: input g0 (A3) @(308,251) /sn:0 /R:3 /w:[ 0 ]
  //: output g12 (S1) @(605,503) /sn:0 /R:3 /w:[ 1 ]

endmodule

module main;    //: root_module
wire w14;    //: /sn:0 {0}(236,9)(275,9)(275,119){1}
wire w4;    //: /sn:0 {0}(312,-61)(327,-61)(327,119){1}
wire w3;    //: /sn:0 {0}(277,-42)(312,-42)(312,119){1}
wire w0;    //: /sn:0 {0}(202,65)(238,65)(238,119){1}
wire w1;    //: /sn:0 {0}(236,38)(257,38)(257,119){1}
wire w8;    //: /sn:0 {0}(202,96)(220,96)(220,119){1}
wire w18;    //: /sn:0 {0}(173,153)(173,159)(208,159){1}
wire w2;    //: /sn:0 {0}(276,-14)(292,-14)(292,119){1}
wire w11;    //: /sn:0 {0}(336,212)(336,249)(353,249)(353,239){1}
wire w12;    //: /sn:0 {0}(285,212)(285,249)(301,249)(301,239){1}
wire w10;    //: /sn:0 {0}(384,212)(384,250)(405,250)(405,240){1}
wire w13;    //: /sn:0 {0}(248,212)(248,248)(260,248)(260,238){1}
wire w5;    //: /sn:0 {0}(312,-90)(345,-90)(345,119){1}
wire w9;    //: /sn:0 {0}(432,98)(442,98)(442,154)(433,154){1}
//: enddecls

  //: switch g8 (w0) @(185,65) /sn:0 /w:[ 0 ] /st:1
  led g4 (.I(w10));   //: @(405,233) /sn:0 /w:[ 1 ] /type:0
  //: switch g13 (w4) @(295,-61) /sn:0 /w:[ 0 ] /st:1
  led g3 (.I(w11));   //: @(353,232) /sn:0 /w:[ 1 ] /type:0
  led g2 (.I(w12));   //: @(301,232) /sn:0 /w:[ 1 ] /type:0
  led g1 (.I(w13));   //: @(260,231) /sn:0 /w:[ 1 ] /type:0
  //: switch g11 (w2) @(259,-14) /sn:0 /w:[ 0 ] /st:1
  //: switch g10 (w14) @(219,9) /sn:0 /w:[ 0 ] /st:1
  //: switch g6 (w9) @(415,98) /sn:0 /w:[ 0 ] /st:0
  //: switch g9 (w1) @(219,38) /sn:0 /w:[ 0 ] /st:1
  //: switch g7 (w8) @(185,96) /sn:0 /w:[ 0 ] /st:1
  //: switch g14 (w5) @(295,-90) /sn:0 /w:[ 0 ] /st:1
  led g5 (.I(w18));   //: @(173,146) /sn:0 /w:[ 0 ] /type:0
  CPA g0 (.B0(w5), .A0(w4), .B1(w3), .A1(w2), .B2(w14), .A2(w1), .B3(w0), .A3(w8), .C0(w9), .C4(w18), .S3(w13), .S2(w12), .S1(w11), .S0(w10));   //: @(209, 120) /sz:(223, 91) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Ti3>1 Ti4>1 Ti5>1 Ti6>1 Ti7>1 Ri0>1 Lo0<1 Bo0<0 Bo1<0 Bo2<0 Bo3<0 ]
  //: switch g12 (w3) @(260,-42) /sn:0 /w:[ 0 ] /st:1

endmodule
