//: version "1.8.7"

module CarryLookahead_Logic(C3, P0, Cout, G0, P3, G1, P1, P2, C2, C1, G3, Cin, G2);
//: interface  /sz:(328, 96) /bd:[ Ti0>G0(286/328) Ti1>P0(267/328) Ti2>G1(210/328) Ti3>P1(189/328) Ti4>G2(139/328) Ti5>P2(117/328) Ti6>G3(55/328) Ti7>P3(28/328) Ri0>Cin(46/96) To0<C3(86/328) To1<C2(159/328) To2<C1(228/328) Lo0<Cout(39/96) ]
input G2;    //: /sn:0 {0}(49,313)(536,313)(536,263)(556,263){1}
input P1;    //: /sn:0 {0}(53,230)(304,230)(304,164)(324,164){1}
output C3;    //: /sn:0 /dp:1 {0}(577,261)(584,261)(584,278)(600,278){1}
//: {2}(604,278)(618,278)(618,269)(622,269){3}
//: {4}(602,280)(602,302)(620,302){5}
input G0;    //: /sn:0 {0}(72,169)(250,169)(250,95)(270,95){1}
output C2;    //: /sn:0 /dp:1 {0}(410,168)(423,168)(423,178)(429,178){1}
//: {2}(433,178)(454,178)(454,177)(456,177){3}
//: {4}(431,180)(431,218)(488,218){5}
input Cin;    //: /sn:0 /dp:1 {0}(200,84)(173,84)(173,65)(85,65){1}
input P3;    //: /sn:0 {0}(40,343)(54,343)(54,307)(620,307){1}
input G1;    //: /sn:0 {0}(51,249)(369,249)(369,170)(389,170){1}
output Cout;    //: /sn:0 /dp:1 {0}(712,334)(742,334)(742,333)(758,333){1}
input G3;    //: /sn:0 {0}(30,372)(681,372)(681,336)(691,336){1}
output C1;    //: /sn:0 /dp:1 {0}(291,93)(303,93)(303,119){1}
//: {2}(305,121)(315,121)(315,159)(324,159){3}
//: {4}(303,123)(303,125)(352,125){5}
input P0;    //: /sn:0 /dp:1 {0}(200,89)(165,89)(165,77)(155,77)(155,145)(72,145){1}
input P2;    //: /sn:0 /dp:1 {0}(488,223)(463,223)(463,272)(453,272)(453,284)(50,284){1}
wire w6;    //: /sn:0 {0}(345,162)(379,162)(379,165)(389,165){1}
wire w3;    //: /sn:0 {0}(509,221)(519,221)(519,258)(556,258){1}
wire w2;    //: /sn:0 {0}(641,305)(651,305)(651,319){1}
//: {2}(653,321)(683,321)(683,331)(691,331){3}
//: {4}(649,321)(625,321){5}
wire w5;    //: /sn:0 {0}(221,87)(260,87)(260,90)(270,90){1}
//: enddecls

  and g8 (.I0(C1), .I1(P1), .Z(w6));   //: @(335,162) /sn:0 /delay:" 1" /w:[ 3 1 0 ]
  or g4 (.I0(w5), .I1(G0), .Z(C1));   //: @(281,93) /sn:0 /delay:" 1" /w:[ 1 1 0 ]
  or g16 (.I0(w3), .I1(G2), .Z(C3));   //: @(567,261) /sn:0 /delay:" 1" /w:[ 1 1 0 ]
  and g3 (.I0(Cin), .I1(P0), .Z(w5));   //: @(211,87) /sn:0 /delay:" 1" /w:[ 0 0 0 ]
  //: output g17 (C3) @(619,269) /sn:0 /w:[ 3 ]
  //: input g2 (P0) @(70,145) /sn:0 /w:[ 1 ]
  //: output g23 (Cout) @(755,333) /sn:0 /w:[ 1 ]
  //: joint g24 (w2) @(651, 321) /w:[ 2 1 4 -1 ]
  //: input g1 (G0) @(70,169) /sn:0 /w:[ 0 ]
  //: input g18 (P3) @(38,343) /sn:0 /w:[ 0 ]
  or g10 (.I0(w6), .I1(G1), .Z(C2));   //: @(400,168) /sn:0 /delay:" 1" /w:[ 1 1 0 ]
  //: input g6 (G1) @(49,249) /sn:0 /w:[ 0 ]
  //: joint g9 (C1) @(303, 121) /w:[ 2 1 -1 4 ]
  //: input g7 (P1) @(51,230) /sn:0 /w:[ 0 ]
  and g22 (.I0(w2), .I1(G3), .Z(Cout));   //: @(702,334) /sn:0 /delay:" 1" /w:[ 3 1 0 ]
  //: input g12 (P2) @(48,284) /sn:0 /w:[ 1 ]
  and g14 (.I0(C2), .I1(P2), .Z(w3));   //: @(499,221) /sn:0 /delay:" 1" /w:[ 5 0 0 ]
  //: output g11 (C2) @(453,177) /sn:0 /w:[ 3 ]
  //: output g5 (C1) @(349,125) /sn:0 /w:[ 5 ]
  //: joint g21 (C3) @(602, 278) /w:[ 2 -1 1 4 ]
  //: input g19 (G3) @(28,372) /sn:0 /w:[ 0 ]
  and g20 (.I0(C3), .I1(P3), .Z(w2));   //: @(631,305) /sn:0 /delay:" 1" /w:[ 5 1 0 ]
  //: joint g15 (C2) @(431, 178) /w:[ 2 -1 1 4 ]
  //: input g0 (Cin) @(83,65) /sn:0 /w:[ 1 ]
  //: input g13 (G2) @(47,313) /sn:0 /w:[ 0 ]

endmodule

module PFA_v1(C, B, P, S, A, G);
//: interface  /sz:(126, 115) /bd:[ Ti0>A(21/126) Ti1>B(82/126) Ri0>C(56/115) Bo0<S(99/126) Bo1<P(11/126) Bo2<G(56/126) ]
input B;    //: /sn:0 {0}(144,200)(161,200){1}
//: {2}(165,200)(202,200)(202,177)(210,177){3}
//: {4}(163,202)(163,320){5}
//: {6}(165,322)(231,322){7}
//: {8}(163,324)(163,361)(240,361){9}
input A;    //: /sn:0 {0}(151,147)(178,147){1}
//: {2}(182,147)(202,147)(202,172)(210,172){3}
//: {4}(180,149)(180,317)(188,317){5}
//: {6}(192,317)(231,317){7}
//: {8}(190,319)(190,356)(240,356){9}
output G;    //: /sn:0 /dp:1 {0}(261,359)(337,359)(337,385)(346,385){1}
input C;    //: /sn:0 {0}(149,271)(266,271)(266,186)(276,186){1}
output P;    //: /sn:0 /dp:1 {0}(252,320)(312,320)(312,319)(322,319){1}
output S;    //: /sn:0 /dp:1 {0}(297,184)(394,184)(394,198)(406,198){1}
wire w2;    //: /sn:0 {0}(231,175)(267,175)(267,181)(276,181){1}
//: enddecls

  xor g4 (.I0(w2), .I1(C), .Z(S));   //: @(287,184) /sn:0 /delay:" 2" /w:[ 1 1 0 ]
  //: joint g8 (B) @(163, 200) /w:[ 2 -1 1 4 ]
  xor g3 (.I0(A), .I1(B), .Z(w2));   //: @(221,175) /sn:0 /delay:" 2" /w:[ 3 3 0 ]
  //: input g2 (C) @(147,271) /sn:0 /w:[ 0 ]
  //: input g1 (B) @(142,200) /sn:0 /w:[ 0 ]
  and g10 (.I0(A), .I1(B), .Z(G));   //: @(251,359) /sn:0 /delay:" 1" /w:[ 9 9 0 ]
  or g6 (.I0(A), .I1(B), .Z(P));   //: @(242,320) /sn:0 /delay:" 1" /w:[ 7 7 0 ]
  //: joint g7 (A) @(180, 147) /w:[ 2 -1 1 4 ]
  //: output g9 (P) @(319,319) /sn:0 /w:[ 1 ]
  //: joint g12 (A) @(190, 317) /w:[ 6 -1 5 8 ]
  //: output g5 (S) @(403,198) /sn:0 /w:[ 1 ]
  //: joint g11 (B) @(163, 322) /w:[ 6 5 -1 8 ]
  //: input g0 (A) @(149,147) /sn:0 /w:[ 0 ]
  //: output g13 (G) @(343,385) /sn:0 /w:[ 1 ]

endmodule

module main;    //: root_module
wire w13;    //: /sn:0 {0}(-477,460)(-477,508){1}
//: {2}(-475,510)(-459,510)(-459,497){3}
//: {4}(-477,512)(-477,519)(-487,519)(-487,559){5}
wire w6;    //: /sn:0 {0}(-276,458)(-276,510)(-335,510)(-335,529){1}
//: {2}(-333,531)(-310,531)(-310,543)(-295,543)(-295,533){3}
//: {4}(-335,533)(-335,559){5}
wire w16;    //: /sn:0 {0}(196,256)(196,322){1}
//: {2}(198,324)(228,324)(228,322){3}
//: {4}(196,326)(196,347)(219,347)(219,355){5}
wire w65;    //: /sn:0 {0}(-1391,442)(-1300,442)(-1300,550){1}
wire w58;    //: /sn:0 {0}(-1582,766)(-1582,598)(-1583,598){1}
//: {2}(-1585,596)(-1585,586)(-1591,586)(-1591,553){3}
//: {4}(-1587,598)(-1602,598){5}
wire w7;    //: /sn:0 {0}(-856,599)(-903,599)(-903,603)(-1013,603){1}
//: {2}(-1017,603)(-1053,603)(-1053,605)(-1061,605){3}
//: {4}(-1015,605)(-1015,813)(-1109,813){5}
wire w88;    //: /sn:0 {0}(-2292,877)(-2292,921)(-2272,921)(-2272,911){1}
wire w50;    //: /sn:0 {0}(-1170,665)(-1170,717)(-1229,717)(-1229,736){1}
//: {2}(-1227,738)(-1204,738)(-1204,750)(-1189,750)(-1189,740){3}
//: {4}(-1229,740)(-1229,766){5}
wire w34;    //: /sn:0 {0}(301,355)(301,327)(334,327)(334,196)(326,196){1}
//: {2}(324,194)(324,184)(323,184)(323,173){3}
//: {4}(322,196)(312,196){5}
wire w81;    //: /sn:0 {0}(-2417,976)(-2417,808)(-2418,808){1}
//: {2}(-2420,806)(-2420,796)(-2426,796)(-2426,763){3}
//: {4}(-2422,808)(-2437,808){5}
wire w59;    //: /sn:0 {0}(-1440,766)(-1440,738)(-1407,738)(-1407,607)(-1415,607){1}
//: {2}(-1417,605)(-1417,595)(-1418,595)(-1418,584){3}
//: {4}(-1419,607)(-1429,607){5}
wire w72;    //: /sn:0 {0}(-1719,476)(-1708,476)(-1708,541){1}
wire w62;    //: /sn:0 {0}(-1189,443)(-1106,443)(-1106,548){1}
wire w39;    //: /sn:0 {0}(-411,559)(-411,524)(-343,524)(-343,402){1}
//: {2}(-343,398)(-343,388)(-349,388)(-349,358){3}
//: {4}(-345,400)(-361,400){5}
wire w4;    //: /sn:0 {0}(571,254)(571,306)(512,306)(512,325){1}
//: {2}(514,327)(537,327)(537,339)(552,339)(552,329){3}
//: {4}(512,329)(512,355){5}
wire w25;    //: /sn:0 {0}(552,72)(574,72)(574,137){1}
wire w56;    //: /sn:0 {0}(-1718,658)(-1718,704){1}
//: {2}(-1716,706)(-1692,706)(-1692,699){3}
//: {4}(-1718,708)(-1718,758)(-1695,758)(-1695,766){5}
wire w82;    //: /sn:0 {0}(-2465,868)(-2465,916)(-2449,916)(-2449,906){1}
wire w36;    //: /sn:0 {0}(-215,606)(-121,606)(-121,398){1}
//: {2}(-119,396)(-30,396)(-30,395)(-9,395){3}
//: {4}(-123,396)(-159,396)(-159,398)(-167,398){5}
wire w3;    //: /sn:0 {0}(609,254)(609,287)(607,287)(607,320){1}
//: {2}(609,322)(675,322)(675,356)(691,356)(691,346){3}
//: {4}(607,324)(607,347)(549,347)(549,355){5}
wire w22;    //: /sn:0 {0}(23,247)(23,293){1}
//: {2}(25,295)(49,295)(49,288){3}
//: {4}(23,297)(23,347)(46,347)(46,355){5}
wire w0;    //: /sn:0 /dp:1 {0}(439,289)(439,299)(458,299)(458,256){1}
wire w60;    //: /sn:0 {0}(-1305,766)(-1305,731)(-1237,731)(-1237,609){1}
//: {2}(-1237,605)(-1237,595)(-1243,595)(-1243,565){3}
//: {4}(-1239,607)(-1255,607){5}
wire w20;    //: /sn:0 {0}(372,67)(380,67)(380,139){1}
wire w71;    //: /sn:0 {0}(-1369,478)(-1361,478)(-1361,550){1}
wire w30;    //: /sn:0 {0}(-824,451)(-824,497){1}
//: {2}(-822,499)(-798,499)(-798,492){3}
//: {4}(-824,501)(-824,551)(-801,551)(-801,559){5}
wire w29;    //: /sn:0 {0}(-779,451)(-779,530){1}
//: {2}(-777,532)(-743,532)(-743,518){3}
//: {4}(-779,534)(-779,551)(-748,551)(-748,559){5}
wire w42;    //: /sn:0 {0}(-601,270)(-580,270)(-580,343){1}
wire w37;    //: /sn:0 {0}(-688,559)(-688,391)(-689,391){1}
//: {2}(-691,389)(-691,379)(-697,379)(-697,346){3}
//: {4}(-693,391)(-708,391){5}
wire w73;    //: /sn:0 {0}(-1630,658)(-1630,706)(-1614,706)(-1614,696){1}
wire w66;    //: /sn:0 {0}(-1556,496)(-1535,496)(-1535,550){1}
wire w12;    //: /sn:0 {0}(-432,460)(-432,503)(-446,503)(-446,538){1}
//: {2}(-444,540)(-438,540)(-438,553)(-423,553)(-423,543){3}
//: {4}(-446,542)(-446,559){5}
wire w18;    //: /sn:0 {0}(185,85)(206,85)(206,139){1}
wire w19;    //: /sn:0 {0}(246,66)(267,66)(267,139){1}
wire w63;    //: /sn:0 {0}(-1302,700)(-1302,710)(-1283,710)(-1283,667){1}
wire w10;    //: /sn:0 {0}(370,256)(370,304){1}
//: {2}(372,306)(388,306)(388,293){3}
//: {4}(370,308)(370,315)(360,315)(360,355){5}
wire w23;    //: /sn:0 {0}(111,247)(111,295)(127,295)(127,285){1}
wire w91;    //: /sn:0 {0}(-1967,875)(-1967,908)(-1969,908)(-1969,941){1}
//: {2}(-1967,943)(-1901,943)(-1901,977)(-1885,977)(-1885,967){3}
//: {4}(-1969,945)(-1969,968)(-2027,968)(-2027,976){5}
wire w84;    //: /sn:0 {0}(-2391,706)(-2370,706)(-2370,760){1}
wire w70;    //: /sn:0 {0}(-1678,393)(-1666,393)(-1666,438)(-1647,438)(-1647,541){1}
wire w54;    //: /sn:0 {0}(-1545,667)(-1545,733){1}
//: {2}(-1543,735)(-1513,735)(-1513,733){3}
//: {4}(-1545,737)(-1545,758)(-1522,758)(-1522,766){5}
wire w86;    //: /sn:0 {0}(-2330,687)(-2309,687)(-2309,760){1}
wire w21;    //: /sn:0 {0}(68,247)(68,326){1}
//: {2}(70,328)(104,328)(104,314){3}
//: {4}(68,330)(68,347)(99,347)(99,355){5}
wire w24;    //: /sn:0 {0}(350,31)(441,31)(441,139){1}
wire w31;    //: /sn:0 {0}(-1132,665)(-1132,698)(-1134,698)(-1134,731){1}
//: {2}(-1132,733)(-1066,733)(-1066,767)(-1050,767)(-1050,757){3}
//: {4}(-1134,735)(-1134,758)(-1192,758)(-1192,766){5}
wire w1;    //: /sn:0 /dp:1 {0}(639,295)(639,305)(652,305)(652,254){1}
wire w68;    //: /sn:0 {0}(-1457,667)(-1457,711)(-1437,711)(-1437,701){1}
wire w32;    //: /sn:0 {0}(632,402)(726,402)(726,194){1}
//: {2}(728,192)(785,192)(785,146)(773,146){3}
//: {4}(724,192)(688,192)(688,194)(680,194){5}
wire w53;    //: /sn:0 {0}(-1500,667)(-1500,708){1}
//: {2}(-1498,710)(-1484,710)(-1484,717)(-1469,717)(-1469,707){3}
//: {4}(-1500,712)(-1500,740)(-1479,740)(-1479,766){5}
wire w46;    //: /sn:0 {0}(-497,235)(-406,235)(-406,343){1}
wire w8;    //: /sn:0 {0}(22,65)(33,65)(33,130){1}
wire w95;    //: /sn:0 {0}(-2024,693)(-2002,693)(-2002,758){1}
wire w89;    //: /sn:0 {0}(-2335,877)(-2335,918){1}
//: {2}(-2333,920)(-2319,920)(-2319,927)(-2304,927)(-2304,917){3}
//: {4}(-2335,922)(-2335,950)(-2314,950)(-2314,976){5}
wire w52;    //: /sn:0 {0}(-1371,667)(-1371,715){1}
//: {2}(-1369,717)(-1353,717)(-1353,704){3}
//: {4}(-1371,719)(-1371,726)(-1381,726)(-1381,766){5}
wire w75;    //: /sn:0 {0}(-2226,652)(-2135,652)(-2135,760){1}
wire w44;    //: /sn:0 {0}(-408,493)(-408,503)(-389,503)(-389,460){1}
wire w27;    //: /sn:0 {0}(-606,460)(-606,501){1}
//: {2}(-604,503)(-590,503)(-590,510)(-575,510)(-575,500){3}
//: {4}(-606,505)(-606,533)(-585,533)(-585,559){5}
wire w17;    //: /sn:0 {0}(284,256)(284,300)(304,300)(304,290){1}
wire w80;    //: /sn:0 {0}(-2513,603)(-2501,603)(-2501,648)(-2482,648)(-2482,751){1}
wire w67;    //: /sn:0 {0}(-1495,477)(-1474,477)(-1474,550){1}
wire w28;    //: /sn:0 {0}(-651,460)(-651,526){1}
//: {2}(-649,528)(-619,528)(-619,526){3}
//: {4}(-651,530)(-651,551)(-628,551)(-628,559){5}
wire w33;    //: /sn:0 {0}(436,355)(436,320)(504,320)(504,198){1}
//: {2}(504,194)(504,184)(498,184)(498,154){3}
//: {4}(502,196)(486,196){5}
wire w35;    //: /sn:0 {0}(159,355)(159,187)(158,187){1}
//: {2}(156,185)(156,175)(150,175)(150,142){3}
//: {4}(154,187)(139,187){5}
wire w69;    //: /sn:0 {0}(-1102,706)(-1102,716)(-1089,716)(-1089,665){1}
wire w49;    //: /sn:0 {0}(-295,236)(-212,236)(-212,341){1}
wire w45;    //: /sn:0 {0}(-475,271)(-467,271)(-467,343){1}
wire w14;    //: /sn:0 {0}(75,27)(94,27)(94,130){1}
wire w78;    //: /sn:0 {0}(-2005,875)(-2005,927)(-2064,927)(-2064,946){1}
//: {2}(-2062,948)(-2039,948)(-2039,960)(-2024,960)(-2024,950){3}
//: {4}(-2064,950)(-2064,976){5}
wire w74;    //: /sn:0 {0}(-2140,976)(-2140,941)(-2072,941)(-2072,819){1}
//: {2}(-2072,815)(-2072,805)(-2078,805)(-2078,775){3}
//: {4}(-2074,817)(-2090,817){5}
wire w2;    //: /sn:0 {0}(-784,186)(-772,186)(-772,231)(-753,231)(-753,334){1}
wire w48;    //: /sn:0 {0}(-295,276)(-273,276)(-273,341){1}
wire w41;    //: /sn:0 {0}(-662,289)(-641,289)(-641,343){1}
wire w11;    //: /sn:0 {0}(-825,269)(-814,269)(-814,334){1}
wire w47;    //: /sn:0 {0}(-208,499)(-208,509)(-195,509)(-195,458){1}
wire w90;    //: /sn:0 {0}(-2204,688)(-2196,688)(-2196,760){1}
wire w85;    //: /sn:0 {0}(-2206,877)(-2206,925){1}
//: {2}(-2204,927)(-2188,927)(-2188,914){3}
//: {4}(-2206,929)(-2206,936)(-2216,936)(-2216,976){5}
wire w83;    //: /sn:0 {0}(-2508,868)(-2508,947){1}
//: {2}(-2506,949)(-2472,949)(-2472,935){3}
//: {4}(-2508,951)(-2508,968)(-2477,968)(-2477,976){5}
wire w15;    //: /sn:0 {0}(241,256)(241,297){1}
//: {2}(243,299)(257,299)(257,306)(272,306)(272,296){3}
//: {4}(241,301)(241,329)(262,329)(262,355){5}
wire w94;    //: /sn:0 {0}(-2618,1006)(-2618,1016)(-2585,1016){1}
wire w92;    //: /sn:0 {0}(-2161,877)(-2161,920)(-2175,920)(-2175,955){1}
//: {2}(-2173,957)(-2167,957)(-2167,970)(-2152,970)(-2152,960){3}
//: {4}(-2175,959)(-2175,976){5}
wire w61;    //: /sn:0 {0}(-1750,806)(-1760,806)(-1760,813)(-1848,813){1}
//: {2}(-1852,813)(-1888,813)(-1888,815)(-1896,815){3}
//: {4}(-1850,815)(-1850,1023)(-1944,1023){5}
wire w55;    //: /sn:0 {0}(-1673,658)(-1673,737){1}
//: {2}(-1671,739)(-1637,739)(-1637,725){3}
//: {4}(-1673,741)(-1673,758)(-1642,758)(-1642,766){5}
wire w38;    //: /sn:0 {0}(-546,559)(-546,531)(-513,531)(-513,400)(-521,400){1}
//: {2}(-523,398)(-523,388)(-524,388)(-524,377){3}
//: {4}(-525,400)(-535,400){5}
wire w5;    //: /sn:0 {0}(-238,458)(-238,491)(-240,491)(-240,524){1}
//: {2}(-238,526)(-172,526)(-172,560)(-156,560)(-156,550){3}
//: {4}(-240,528)(-240,551)(-298,551)(-298,559){5}
wire w87;    //: /sn:0 {0}(-2275,976)(-2275,948)(-2242,948)(-2242,817)(-2250,817){1}
//: {2}(-2252,815)(-2252,805)(-2253,805)(-2253,794){3}
//: {4}(-2254,817)(-2264,817){5}
wire w64;    //: /sn:0 {0}(-1189,483)(-1167,483)(-1167,548){1}
wire w43;    //: /sn:0 {0}(-563,460)(-563,504)(-543,504)(-543,494){1}
wire w97;    //: /sn:0 {0}(-2137,910)(-2137,920)(-2118,920)(-2118,877){1}
wire w96;    //: /sn:0 {0}(-1937,916)(-1937,926)(-1924,926)(-1924,875){1}
wire w76;    //: /sn:0 {0}(-2380,877)(-2380,943){1}
//: {2}(-2378,945)(-2348,945)(-2348,943){3}
//: {4}(-2380,947)(-2380,968)(-2357,968)(-2357,976){5}
wire w9;    //: /sn:0 {0}(415,256)(415,299)(401,299)(401,334){1}
//: {2}(403,336)(409,336)(409,349)(424,349)(424,339){3}
//: {4}(401,338)(401,355){5}
wire w26;    //: /sn:0 {0}(552,32)(635,32)(635,137){1}
wire w79;    //: /sn:0 {0}(-2554,686)(-2543,686)(-2543,751){1}
wire w77;    //: /sn:0 {0}(-2024,653)(-1941,653)(-1941,758){1}
wire w57;    //: /sn:0 {0}(-2553,868)(-2553,914){1}
//: {2}(-2551,916)(-2527,916)(-2527,909){3}
//: {4}(-2553,918)(-2553,968)(-2530,968)(-2530,976){5}
wire w51;    //: /sn:0 {0}(-1326,667)(-1326,710)(-1340,710)(-1340,745){1}
//: {2}(-1338,747)(-1332,747)(-1332,760)(-1317,760)(-1317,750){3}
//: {4}(-1340,749)(-1340,766){5}
wire w40;    //: /sn:0 {0}(-736,451)(-736,499)(-720,499)(-720,489){1}
//: enddecls

  //: switch g8 (w8) @(5,65) /sn:0 /w:[ 0 ] /st:0
  CarryLookahead_Logic g4 (.G0(w3), .P0(w4), .G1(w9), .P1(w10), .G2(w15), .P2(w16), .G3(w21), .P3(w22), .Cin(w32), .C3(w35), .C2(w34), .C1(w33), .Cout(w36));   //: @(-8, 356) /sz:(639, 96) /sn:0 /p:[ Ti0>5 Ti1>5 Ti2>5 Ti3>5 Ti4>5 Ti5>5 Ti6>5 Ti7>5 Ri0>0 To0<0 To1<0 To2<0 Lo0<3 ]
  led g116 (.I(w60));   //: @(-1243,558) /sn:0 /w:[ 3 ] /type:0
  //: switch g157 (w95) @(-2041,693) /sn:0 /w:[ 0 ] /st:1
  //: joint g17 (w33) @(504, 196) /w:[ -1 2 4 1 ]
  //: joint g137 (w81) @(-2420, 808) /w:[ 1 2 4 -1 ]
  led g30 (.I(w9));   //: @(424,332) /sn:0 /w:[ 3 ] /type:0
  //: joint g74 (w38) @(-523, 400) /w:[ 1 2 4 -1 ]
  led g92 (.I(w54));   //: @(-1513,726) /sn:0 /w:[ 3 ] /type:0
  PFA_v1 g130 (.A(w79), .B(w80), .C(w81), .S(w82), .P(w57), .G(w83));   //: @(-2564, 752) /sz:(126, 115) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>5 Bo0<0 Bo1<0 Bo2<0 ]
  PFA_v1 g1 (.A(w20), .B(w24), .C(w33), .S(w0), .P(w10), .G(w9));   //: @(359, 140) /sz:(126, 115) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>5 Bo0<1 Bo1<0 Bo2<0 ]
  //: switch g77 (w49) @(-312,236) /sn:0 /w:[ 0 ] /st:0
  PFA_v1 g111 (.A(w72), .B(w70), .C(w58), .S(w73), .P(w56), .G(w55));   //: @(-1729, 542) /sz:(126, 115) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>5 Bo0<0 Bo1<0 Bo2<0 ]
  //: joint g144 (w83) @(-2508, 949) /w:[ 2 1 -1 4 ]
  led g51 (.I(w44));   //: @(-408,486) /sn:0 /w:[ 0 ] /type:0
  //: joint g161 (w91) @(-1969, 943) /w:[ 2 1 -1 4 ]
  //: switch g70 (w48) @(-312,276) /sn:0 /w:[ 0 ] /st:1
  led g149 (.I(w88));   //: @(-2272,904) /sn:0 /w:[ 1 ] /type:0
  led g25 (.I(w1));   //: @(639,288) /sn:0 /w:[ 0 ] /type:0
  //: switch g10 (w18) @(168,85) /sn:0 /w:[ 0 ] /st:0
  //: joint g65 (w30) @(-824, 499) /w:[ 2 1 -1 4 ]
  //: joint g103 (w60) @(-1237, 607) /w:[ -1 2 4 1 ]
  led g64 (.I(w28));   //: @(-619,519) /sn:0 /w:[ 3 ] /type:0
  PFA_v1 g49 (.A(w41), .B(w42), .C(w38), .S(w43), .P(w28), .G(w27));   //: @(-662, 344) /sz:(126, 115) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>5 Bo0<0 Bo1<0 Bo2<0 ]
  led g72 (.I(w58));   //: @(-1591,546) /sn:0 /w:[ 3 ] /type:0
  CarryLookahead_Logic g142 (.G0(w91), .P0(w78), .G1(w92), .P1(w85), .G2(w89), .P2(w76), .G3(w83), .P3(w57), .Cin(w61), .C3(w81), .C2(w87), .C1(w74), .Cout(w94));   //: @(-2584, 977) /sz:(639, 96) /sn:0 /p:[ Ti0>5 Ti1>5 Ti2>5 Ti3>5 Ti4>5 Ti5>5 Ti6>5 Ti7>5 Ri0>5 To0<0 To1<0 To2<0 Lo0<1 ]
  led g136 (.I(w81));   //: @(-2426,756) /sn:0 /w:[ 3 ] /type:0
  //: joint g6 (w32) @(726, 192) /w:[ 2 -1 4 1 ]
  //: joint g35 (w15) @(241, 299) /w:[ 2 1 -1 4 ]
  led g56 (.I(w47));   //: @(-208,492) /sn:0 /w:[ 0 ] /type:0
  //: joint g58 (w36) @(-121, 396) /w:[ 2 -1 4 1 ]
  //: switch g7 (w2) @(-801,186) /sn:0 /w:[ 0 ] /st:0
  led g124 (.I(w57));   //: @(-2527,902) /sn:0 /w:[ 3 ] /type:0
  //: joint g98 (w58) @(-1585, 598) /w:[ 1 2 4 -1 ]
  //: switch g67 (w45) @(-492,271) /sn:0 /w:[ 0 ] /st:1
  //: joint g85 (w59) @(-1417, 607) /w:[ 1 2 4 -1 ]
  led g126 (.I(w76));   //: @(-2348,936) /sn:0 /w:[ 3 ] /type:0
  //: joint g33 (w10) @(370, 306) /w:[ 2 1 -1 4 ]
  //: joint g54 (w6) @(-335, 531) /w:[ 2 1 -1 4 ]
  led g40 (.I(w22));   //: @(49,281) /sn:0 /w:[ 3 ] /type:0
  //: joint g52 (w29) @(-779, 532) /w:[ 2 1 -1 4 ]
  //: joint g81 (w28) @(-651, 528) /w:[ 2 1 -1 4 ]
  PFA_v1 g163 (.A(w90), .B(w75), .C(w74), .S(w97), .P(w85), .G(w92));   //: @(-2217, 761) /sz:(126, 115) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>5 Bo0<1 Bo1<0 Bo2<0 ]
  //: joint g132 (w74) @(-2072, 817) /w:[ -1 2 4 1 ]
  //: switch g12 (w20) @(355,67) /sn:0 /w:[ 0 ] /st:1
  //: joint g108 (w54) @(-1545, 735) /w:[ 2 1 -1 4 ]
  led g131 (.I(w85));   //: @(-2188,907) /sn:0 /w:[ 3 ] /type:0
  //: joint g106 (w55) @(-1673, 739) /w:[ 2 1 -1 4 ]
  //: joint g96 (w7) @(-1015, 603) /w:[ 1 -1 2 4 ]
  //: joint g19 (w34) @(324, 196) /w:[ 1 2 4 -1 ]
  PFA_v1 g114 (.A(w64), .B(w62), .C(w7), .S(w69), .P(w50), .G(w31));   //: @(-1188, 549) /sz:(126, 115) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>3 Bo0<1 Bo1<0 Bo2<0 ]
  led g117 (.I(w68));   //: @(-1437,694) /sn:0 /w:[ 1 ] /type:0
  led g78 (.I(w29));   //: @(-743,511) /sn:0 /w:[ 3 ] /type:0
  //: joint g125 (w57) @(-2553, 916) /w:[ 2 1 -1 4 ]
  //: switch g155 (w79) @(-2571,686) /sn:0 /w:[ 0 ] /st:0
  //: joint g63 (w13) @(-477, 510) /w:[ 2 1 -1 4 ]
  led g93 (.I(w51));   //: @(-1317,743) /sn:0 /w:[ 3 ] /type:0
  //: switch g105 (w72) @(-1736,476) /sn:0 /w:[ 0 ] /st:0
  led g113 (.I(w55));   //: @(-1637,718) /sn:0 /w:[ 3 ] /type:0
  PFA_v1 g0 (.A(w25), .B(w26), .C(w32), .S(w1), .P(w4), .G(w3));   //: @(553, 138) /sz:(126, 115) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>5 Bo0<1 Bo1<0 Bo2<0 ]
  led g38 (.I(w21));   //: @(104,307) /sn:0 /w:[ 3 ] /type:0
  led g43 (.I(w39));   //: @(-349,351) /sn:0 /w:[ 3 ] /type:0
  //: switch g101 (w67) @(-1512,477) /sn:0 /w:[ 0 ] /st:1
  led g48 (.I(w43));   //: @(-543,487) /sn:0 /w:[ 1 ] /type:0
  //: joint g37 (w16) @(196, 324) /w:[ 2 1 -1 4 ]
  //: joint g80 (w5) @(-240, 526) /w:[ 2 1 -1 4 ]
  led g95 (.I(w69));   //: @(-1102,699) /sn:0 /w:[ 0 ] /type:0
  //: joint g120 (w31) @(-1134, 733) /w:[ 2 1 -1 4 ]
  PFA_v1 g122 (.A(w71), .B(w65), .C(w60), .S(w63), .P(w52), .G(w51));   //: @(-1382, 551) /sz:(126, 115) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>5 Bo0<1 Bo1<0 Bo2<0 ]
  led g76 (.I(w13));   //: @(-459,490) /sn:0 /w:[ 3 ] /type:0
  led g152 (.I(w92));   //: @(-2152,953) /sn:0 /w:[ 3 ] /type:0
  CarryLookahead_Logic g44 (.G0(w5), .P0(w6), .G1(w12), .P1(w13), .G2(w27), .P2(w28), .G3(w29), .P3(w30), .Cin(w36), .C3(w37), .C2(w38), .C1(w39), .Cout(w7));   //: @(-855, 560) /sz:(639, 96) /sn:0 /p:[ Ti0>5 Ti1>5 Ti2>5 Ti3>5 Ti4>5 Ti5>5 Ti6>5 Ti7>5 Ri0>0 To0<0 To1<0 To2<0 Lo0<0 ]
  led g75 (.I(w37));   //: @(-697,339) /sn:0 /w:[ 3 ] /type:0
  led g159 (.I(w97));   //: @(-2137,903) /sn:0 /w:[ 0 ] /type:0
  led g16 (.I(w33));   //: @(498,147) /sn:0 /w:[ 3 ] /type:0
  PFA_v1 g3 (.A(w8), .B(w14), .C(w35), .S(w23), .P(w22), .G(w21));   //: @(12, 131) /sz:(126, 115) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>5 Bo0<0 Bo1<0 Bo2<0 ]
  led g47 (.I(w5));   //: @(-156,543) /sn:0 /w:[ 3 ] /type:0
  //: joint g143 (w76) @(-2380, 945) /w:[ 2 1 -1 4 ]
  led g26 (.I(w3));   //: @(691,339) /sn:0 /w:[ 3 ] /type:0
  //: switch g90 (w65) @(-1408,442) /sn:0 /w:[ 0 ] /st:0
  led g109 (.I(w56));   //: @(-1692,692) /sn:0 /w:[ 3 ] /type:0
  //: switch g158 (w86) @(-2347,687) /sn:0 /w:[ 0 ] /st:1
  PFA_v1 g2 (.A(w18), .B(w19), .C(w34), .S(w17), .P(w16), .G(w15));   //: @(185, 140) /sz:(126, 115) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>5 Bo0<0 Bo1<0 Bo2<0 ]
  //: joint g128 (w78) @(-2064, 948) /w:[ 2 1 -1 4 ]
  led g23 (.I(w17));   //: @(304,283) /sn:0 /w:[ 1 ] /type:0
  //: joint g91 (w56) @(-1718, 706) /w:[ 2 1 -1 4 ]
  //: switch g141 (w80) @(-2530,603) /sn:0 /w:[ 0 ] /st:0
  led g24 (.I(w0));   //: @(439,282) /sn:0 /w:[ 0 ] /type:0
  //: joint g39 (w21) @(68, 328) /w:[ 2 1 -1 4 ]
  //: switch g86 (w62) @(-1206,443) /sn:0 /w:[ 0 ] /st:0
  //: joint g104 (w50) @(-1229, 738) /w:[ 2 1 -1 4 ]
  //: switch g127 (w77) @(-2041,653) /sn:0 /w:[ 0 ] /st:0
  //: joint g29 (w4) @(512, 327) /w:[ 2 1 -1 4 ]
  //: joint g60 (w27) @(-606, 503) /w:[ 2 1 -1 4 ]
  //: switch g110 (w66) @(-1573,496) /sn:0 /w:[ 0 ] /st:0
  led g121 (.I(w52));   //: @(-1353,697) /sn:0 /w:[ 3 ] /type:0
  led g18 (.I(w34));   //: @(323,166) /sn:0 /w:[ 3 ] /type:0
  //: switch g82 (w46) @(-514,235) /sn:0 /w:[ 0 ] /st:0
  PFA_v1 g94 (.A(w66), .B(w67), .C(w59), .S(w68), .P(w54), .G(w53));   //: @(-1556, 551) /sz:(126, 115) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>5 Bo0<0 Bo1<0 Bo2<0 ]
  led g119 (.I(w59));   //: @(-1418,577) /sn:0 /w:[ 3 ] /type:0
  led g154 (.I(w94));   //: @(-2618,999) /sn:0 /w:[ 0 ] /type:0
  led g107 (.I(w53));   //: @(-1469,700) /sn:0 /w:[ 3 ] /type:0
  led g50 (.I(w12));   //: @(-423,536) /sn:0 /w:[ 3 ] /type:0
  PFA_v1 g133 (.A(w84), .B(w86), .C(w87), .S(w88), .P(w76), .G(w89));   //: @(-2391, 761) /sz:(126, 115) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>5 Bo0<0 Bo1<0 Bo2<0 ]
  //: switch g9 (w14) @(58,27) /sn:0 /w:[ 0 ] /st:0
  led g68 (.I(w6));   //: @(-295,526) /sn:0 /w:[ 3 ] /type:0
  //: joint g73 (w37) @(-691, 391) /w:[ 1 2 4 -1 ]
  led g22 (.I(w23));   //: @(127,278) /sn:0 /w:[ 1 ] /type:0
  //: joint g31 (w9) @(401, 336) /w:[ 2 1 -1 4 ]
  //: switch g71 (w42) @(-618,270) /sn:0 /w:[ 0 ] /st:1
  //: switch g102 (w71) @(-1386,478) /sn:0 /w:[ 0 ] /st:1
  led g59 (.I(w74));   //: @(-2078,768) /sn:0 /w:[ 3 ] /type:0
  //: joint g87 (w53) @(-1500, 710) /w:[ 2 1 -1 4 ]
  CarryLookahead_Logic g83 (.G0(w31), .P0(w50), .G1(w51), .P1(w52), .G2(w53), .P2(w54), .G3(w55), .P3(w56), .Cin(w7), .C3(w58), .C2(w59), .C1(w60), .Cout(w61));   //: @(-1749, 767) /sz:(639, 96) /sn:0 /p:[ Ti0>5 Ti1>5 Ti2>5 Ti3>5 Ti4>5 Ti5>5 Ti6>5 Ti7>5 Ri0>5 To0<0 To1<0 To2<0 Lo0<0 ]
  //: switch g99 (w70) @(-1695,393) /sn:0 /w:[ 0 ] /st:0
  led g36 (.I(w16));   //: @(228,315) /sn:0 /w:[ 3 ] /type:0
  //: joint g41 (w22) @(23, 295) /w:[ 2 1 -1 4 ]
  //: joint g45 (w39) @(-343, 400) /w:[ -1 2 4 1 ]
  led g156 (.I(w83));   //: @(-2472,928) /sn:0 /w:[ 3 ] /type:0
  //: switch g138 (w90) @(-2221,688) /sn:0 /w:[ 0 ] /st:1
  //: switch g42 (w11) @(-842,269) /sn:0 /w:[ 0 ] /st:0
  led g69 (.I(w27));   //: @(-575,493) /sn:0 /w:[ 3 ] /type:0
  //: joint g151 (w85) @(-2206, 927) /w:[ 2 1 -1 4 ]
  led g66 (.I(w30));   //: @(-798,485) /sn:0 /w:[ 3 ] /type:0
  led g153 (.I(w78));   //: @(-2024,943) /sn:0 /w:[ 3 ] /type:0
  //: joint g146 (w92) @(-2175, 957) /w:[ 2 1 -1 4 ]
  led g28 (.I(w4));   //: @(552,322) /sn:0 /w:[ 3 ] /type:0
  led g34 (.I(w15));   //: @(272,289) /sn:0 /w:[ 3 ] /type:0
  PFA_v1 g46 (.A(w11), .B(w2), .C(w37), .S(w40), .P(w30), .G(w29));   //: @(-835, 335) /sz:(126, 115) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>5 Bo0<0 Bo1<0 Bo2<0 ]
  //: switch g57 (w41) @(-679,289) /sn:0 /w:[ 0 ] /st:0
  PFA_v1 g150 (.A(w95), .B(w77), .C(w61), .S(w96), .P(w78), .G(w91));   //: @(-2023, 759) /sz:(126, 115) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>3 Bo0<1 Bo1<0 Bo2<0 ]
  //: switch g14 (w25) @(535,72) /sn:0 /w:[ 0 ] /st:1
  //: switch g11 (w19) @(229,66) /sn:0 /w:[ 0 ] /st:1
  //: switch g5 (w32) @(756,146) /sn:0 /w:[ 3 ] /st:0
  led g84 (.I(w31));   //: @(-1050,750) /sn:0 /w:[ 3 ] /type:0
  //: joint g118 (w51) @(-1340, 747) /w:[ 2 1 -1 4 ]
  led g112 (.I(w73));   //: @(-1614,689) /sn:0 /w:[ 1 ] /type:0
  //: joint g21 (w35) @(156, 187) /w:[ 1 2 4 -1 ]
  led g61 (.I(w40));   //: @(-720,482) /sn:0 /w:[ 1 ] /type:0
  //: switch g123 (w75) @(-2243,652) /sn:0 /w:[ 0 ] /st:0
  led g20 (.I(w35));   //: @(150,135) /sn:0 /w:[ 3 ] /type:0
  led g32 (.I(w10));   //: @(388,286) /sn:0 /w:[ 3 ] /type:0
  PFA_v1 g79 (.A(w48), .B(w49), .C(w36), .S(w47), .P(w6), .G(w5));   //: @(-294, 342) /sz:(126, 115) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>5 Bo0<1 Bo1<0 Bo2<0 ]
  //: joint g115 (w52) @(-1371, 717) /w:[ 2 1 -1 4 ]
  led g145 (.I(w91));   //: @(-1885,960) /sn:0 /w:[ 3 ] /type:0
  led g134 (.I(w87));   //: @(-2253,787) /sn:0 /w:[ 3 ] /type:0
  led g97 (.I(w50));   //: @(-1189,733) /sn:0 /w:[ 3 ] /type:0
  led g148 (.I(w82));   //: @(-2449,899) /sn:0 /w:[ 1 ] /type:0
  //: switch g129 (w84) @(-2408,706) /sn:0 /w:[ 0 ] /st:0
  //: switch g15 (w26) @(535,32) /sn:0 /w:[ 0 ] /st:0
  //: switch g89 (w64) @(-1206,483) /sn:0 /w:[ 0 ] /st:1
  //: joint g147 (w61) @(-1850, 813) /w:[ 1 -1 2 4 ]
  //: joint g27 (w3) @(607, 322) /w:[ 2 1 -1 4 ]
  led g160 (.I(w96));   //: @(-1937,909) /sn:0 /w:[ 0 ] /type:0
  //: joint g62 (w12) @(-446, 540) /w:[ 2 1 -1 4 ]
  led g55 (.I(w38));   //: @(-524,370) /sn:0 /w:[ 3 ] /type:0
  led g88 (.I(w63));   //: @(-1302,693) /sn:0 /w:[ 0 ] /type:0
  //: joint g140 (w89) @(-2335, 920) /w:[ 2 1 -1 4 ]
  //: joint g139 (w87) @(-2252, 817) /w:[ 1 2 4 -1 ]
  led g135 (.I(w89));   //: @(-2304,910) /sn:0 /w:[ 3 ] /type:0
  //: switch g13 (w24) @(333,31) /sn:0 /w:[ 0 ] /st:0
  PFA_v1 g53 (.A(w45), .B(w46), .C(w39), .S(w44), .P(w13), .G(w12));   //: @(-488, 344) /sz:(126, 115) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>5 Bo0<1 Bo1<0 Bo2<0 ]

endmodule
