//: version "1.8.7"

module ha(S, CO, B, A);
//: interface  /sz:(55, 65) /bd:[ Li0>A(20/65) Li1>B(35/65) Ro0<S(21/65) Ro1<CO(41/65) ]
input B;    //: /sn:0 {0}(170,290)(233,290)(233,291)(292,291){1}
//: {2}(296,291)(373,291)(373,258)(377,258){3}
//: {4}(294,289)(294,259)(302,259){5}
input A;    //: /sn:0 {0}(171,218)(275,218){1}
//: {2}(279,218)(365,218)(365,253)(377,253){3}
//: {4}(277,220)(277,254)(302,254){5}
output CO;    //: /sn:0 /dp:1 {0}(323,257)(352,257){1}
output S;    //: /sn:0 {0}(428,255)(407,255)(407,256)(398,256){1}
//: enddecls

  xor g4 (.I0(A), .I1(B), .Z(S));   //: @(388,256) /sn:0 /delay:" 2" /w:[ 3 3 1 ]
  //: output g3 (S) @(425,255) /sn:0 /w:[ 0 ]
  //: output g2 (CO) @(349,257) /sn:0 /w:[ 1 ]
  //: input g1 (B) @(168,290) /sn:0 /w:[ 0 ]
  //: joint g6 (A) @(277, 218) /w:[ 2 -1 1 4 ]
  //: joint g7 (B) @(294, 291) /w:[ 2 4 1 -1 ]
  and g5 (.I0(A), .I1(B), .Z(CO));   //: @(313,257) /sn:0 /tech:unit /w:[ 5 5 0 ]
  //: input g0 (A) @(169,218) /sn:0 /w:[ 0 ]

endmodule

module RCA_4b(Y0, Z0, X3, X2, X1, Z2, Y2, Y3, Z1, Z4, Y1, Z3, Z6, X0, Z7, Z5);
//: interface  /sz:(128, 136) /bd:[ Ti0>Y3(14/128) Ti1>Y2(25/128) Ti2>Y1(34/128) Ti3>Y0(47/128) Ti4>X3(87/128) Ti5>X2(98/128) Ti6>X1(107/128) Ti7>X0(116/128) Bo0<Z7(41/128) Bo1<Z6(51/128) Bo2<Z5(60/128) Bo3<Z4(70/128) Bo4<Z3(81/128) Bo5<Z2(92/128) Bo6<Z1(104/128) Bo7<Z0(116/128) ]
input X1;    //: /sn:0 /dp:1 {0}(335,159)(335,123){1}
//: {2}(335,119)(335,79){3}
//: {4}(333,121)(293,121)(293,226){5}
input Y3;    //: /sn:0 {0}(545,334)(535,334){1}
input Y2;    //: /sn:0 {0}(548,269)(538,269){1}
output Z0;    //: /sn:0 /dp:1 {0}(426,177)(426,473){1}
output Z3;    //: /sn:0 /dp:1 {0}(296,476)(296,486){1}
input X2;    //: /sn:0 /dp:1 {0}(252,159)(252,124){1}
//: {2}(252,120)(252,80){3}
//: {4}(250,122)(204,122)(204,224){5}
output Z4;    //: /sn:0 /dp:1 {0}(242,475)(242,485){1}
output Z6;    //: /sn:0 /dp:1 {0}(133,495)(133,505){1}
output Z5;    //: /sn:0 /dp:1 {0}(182,489)(182,499){1}
input X0;    //: /sn:0 {0}(424,78)(424,120){1}
//: {2}(422,122)(377,122)(377,224){3}
//: {4}(424,124)(424,156){5}
output Z7;    //: /sn:0 /dp:1 {0}(99,501)(99,511){1}
output Z2;    //: /sn:0 /dp:1 {0}(350,470)(350,480){1}
output Z1;    //: /sn:0 /dp:1 {0}(378,351)(378,476){1}
input Y0;    //: /sn:0 {0}(544,146)(431,146){1}
//: {2}(427,146)(342,146){3}
//: {4}(338,146)(259,146){5}
//: {6}(255,146)(176,146)(176,160){7}
//: {8}(257,148)(257,159){9}
//: {10}(340,148)(340,159){11}
//: {12}(429,148)(429,156){13}
input X3;    //: /sn:0 /dp:1 {0}(171,160)(171,126){1}
//: {2}(171,122)(171,80){3}
//: {4}(169,124)(128,124)(128,224){5}
input Y1;    //: /sn:0 /dp:1 {0}(382,224)(382,217){1}
//: {2}(384,215)(546,215){3}
//: {4}(380,215)(300,215){5}
//: {6}(296,215)(211,215){7}
//: {8}(209,213)(209,224){9}
//: {10}(207,215)(133,215)(133,224){11}
//: {12}(298,217)(298,226){13}
wire w13;    //: /sn:0 {0}(128,354)(128,364){1}
wire w6;    //: /sn:0 {0}(337,180)(337,284)(364,284)(364,294){1}
wire w7;    //: /sn:0 {0}(379,245)(379,294){1}
wire w4;    //: /sn:0 {0}(256,328)(226,328){1}
wire w3;    //: /sn:0 {0}(356,351)(356,360)(326,360)(326,324)(302,324){1}
wire w18;    //: /sn:0 {0}(130,245)(130,279)(113,279)(113,311){1}
wire w12;    //: /sn:0 {0}(173,181)(173,299)(178,299)(178,309){1}
wire w10;    //: /sn:0 {0}(198,351)(198,361){1}
wire w8;    //: /sn:0 {0}(169,330)(153,330)(153,301)(123,301)(123,311){1}
wire w2;    //: /sn:0 {0}(113,354)(113,364){1}
wire w11;    //: /sn:0 {0}(295,247)(295,294)(289,294)(289,304){1}
wire w15;    //: /sn:0 {0}(206,245)(206,299)(210,299)(210,309){1}
wire w5;    //: /sn:0 {0}(278,349)(278,359){1}
wire w9;    //: /sn:0 {0}(254,180)(254,294)(264,294)(264,304){1}
//: enddecls

  //: input g4 (Y0) @(546,146) /sn:0 /R:2 /w:[ 0 ]
  //: output g8 (Z0) @(426,470) /sn:0 /R:3 /w:[ 1 ]
  //: input g3 (X3) @(171,78) /sn:0 /R:3 /w:[ 3 ]
  and g16 (.I0(Y0), .I1(X0), .Z(Z0));   //: @(426,167) /sn:0 /R:3 /w:[ 13 5 0 ]
  and g26 (.I0(Y1), .I1(X2), .Z(w15));   //: @(206,235) /sn:0 /R:3 /w:[ 9 5 0 ]
  ha g17 (.B(w6), .A(w7), .CO(w3), .S(Z1));   //: @(335, 295) /sz:(65, 55) /sn:0 /p:[ Ti0>1 Ti1>1 Bo0<0 Bo1<0 ]
  //: input g2 (X2) @(252,78) /sn:0 /R:3 /w:[ 3 ]
  //: joint g30 (Y1) @(209, 215) /w:[ 7 8 10 -1 ]
  //: joint g23 (Y0) @(257, 146) /w:[ 5 -1 6 8 ]
  and g24 (.I0(Y1), .I1(X0), .Z(w7));   //: @(379,235) /sn:0 /R:3 /w:[ 0 3 0 ]
  //: input g1 (X1) @(335,77) /sn:0 /R:3 /w:[ 3 ]
  //: joint g29 (Y1) @(298, 215) /w:[ 5 -1 6 12 ]
  and g18 (.I0(Y0), .I1(X1), .Z(w6));   //: @(337,170) /sn:0 /R:3 /w:[ 11 0 0 ]
  and g25 (.I0(Y1), .I1(X1), .Z(w11));   //: @(295,237) /sn:0 /R:3 /w:[ 13 5 0 ]
  //: output g10 (Z2) @(350,477) /sn:0 /R:3 /w:[ 1 ]
  //: input g6 (Y2) @(550,269) /sn:0 /R:2 /w:[ 0 ]
  FA g35 (.A(w9), .B(w11), .Cin(w3), .Cout(w4), .S(w5));   //: @(257, 305) /sz:(44, 43) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  //: input g7 (Y3) @(547,334) /sn:0 /R:2 /w:[ 0 ]
  //: output g9 (Z1) @(378,473) /sn:0 /R:3 /w:[ 1 ]
  //: joint g31 (X3) @(171, 124) /w:[ -1 2 4 1 ]
  //: joint g22 (Y0) @(340, 146) /w:[ 3 -1 4 10 ]
  FA g36 (.A(w12), .B(w15), .Cin(w4), .Cout(w8), .S(w10));   //: @(170, 310) /sz:(55, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  //: joint g33 (X1) @(335, 121) /w:[ -1 2 4 1 ]
  //: output g12 (Z4) @(242,482) /sn:0 /R:3 /w:[ 1 ]
  //: joint g34 (X0) @(424, 122) /w:[ -1 1 2 4 ]
  //: joint g28 (Y1) @(382, 215) /w:[ 2 -1 4 1 ]
  //: input g5 (Y1) @(548,215) /sn:0 /R:2 /w:[ 3 ]
  //: output g11 (Z3) @(296,483) /sn:0 /R:3 /w:[ 1 ]
  //: output g14 (Z6) @(133,502) /sn:0 /R:3 /w:[ 1 ]
  //: joint g21 (Y0) @(429, 146) /w:[ 1 -1 2 12 ]
  and g19 (.I0(Y0), .I1(X2), .Z(w9));   //: @(254,170) /sn:0 /R:3 /w:[ 9 0 0 ]
  //: joint g32 (X2) @(252, 122) /w:[ -1 2 4 1 ]
  and g20 (.I0(Y0), .I1(X3), .Z(w12));   //: @(173,171) /sn:0 /R:3 /w:[ 7 0 0 ]
  //: input g0 (X0) @(424,76) /sn:0 /R:3 /w:[ 0 ]
  //: output g15 (Z7) @(99,508) /sn:0 /R:3 /w:[ 1 ]
  and g27 (.I0(Y1), .I1(X3), .Z(w18));   //: @(130,235) /sn:0 /R:3 /w:[ 11 5 0 ]
  ha g37 (.B(w8), .A(w18), .CO(w13), .S(w2));   //: @(99, 312) /sz:(46, 41) /sn:0 /p:[ Ti0>1 Ti1>1 Bo0<0 Bo1<0 ]
  //: output g13 (Z5) @(182,496) /sn:0 /R:3 /w:[ 1 ]

endmodule

module main;    //: root_module
wire w6;    //: /sn:0 {0}(180,118)(180,128){1}
wire w13;    //: /sn:0 {0}(215,276)(215,266){1}
wire w7;    //: /sn:0 {0}(169,117)(169,128){1}
wire w4;    //: /sn:0 {0}(202,118)(202,128){1}
wire w0;    //: /sn:0 {0}(271,118)(271,128){1}
wire w3;    //: /sn:0 {0}(242,118)(242,128){1}
wire w12;    //: /sn:0 {0}(225,276)(225,266){1}
wire w10;    //: /sn:0 {0}(247,276)(247,266){1}
wire w1;    //: /sn:0 {0}(262,118)(262,128){1}
wire w8;    //: /sn:0 {0}(271,276)(271,266){1}
wire w14;    //: /sn:0 {0}(206,276)(206,266){1}
wire w2;    //: /sn:0 {0}(253,118)(253,128){1}
wire w11;    //: /sn:0 {0}(236,276)(236,266){1}
wire w15;    //: /sn:0 {0}(196,276)(196,266){1}
wire w5;    //: /sn:0 {0}(189,118)(189,128){1}
wire w9;    //: /sn:0 {0}(259,276)(259,266){1}
//: enddecls

  RCA_4b g0 (.Y3(w7), .Y2(w6), .Y1(w5), .Y0(w4), .X3(w3), .X2(w2), .X1(w1), .X0(w0), .Z7(w15), .Z6(w14), .Z5(w13), .Z4(w12), .Z3(w11), .Z2(w10), .Z1(w9), .Z0(w8));   //: @(155, 129) /sz:(128, 136) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Ti3>1 Ti4>1 Ti5>1 Ti6>1 Ti7>1 Bo0<1 Bo1<1 Bo2<1 Bo3<1 Bo4<1 Bo5<1 Bo6<1 Bo7<1 ]

endmodule

module FA(Cout, S, Cin, B, A);
//: interface  /sz:(225, 114) /bd:[ Ti0>B(166/225) Ti1>A(36/225) Ri0>Cin(52/114) Lo0<Cout(58/114) Bo0<S(117/225) ]
input B;    //: /sn:0 {0}(143,173)(159,173){1}
//: {2}(163,173)(176,173)(176,104)(186,104){3}
//: {4}(161,175)(161,176)(242,176)(242,152)(252,152){5}
input A;    //: /sn:0 {0}(130,98)(150,98){1}
//: {2}(154,98)(176,98)(176,99)(186,99){3}
//: {4}(152,100)(152,147)(252,147){5}
input Cin;    //: /sn:0 {0}(143,199)(213,199)(213,125){1}
//: {2}(215,123)(225,123)(225,124)(253,124){3}
//: {4}(213,121)(213,107)(223,107){5}
output Cout;    //: /sn:0 /dp:1 {0}(324,137)(347,137)(347,136)(357,136){1}
output S;    //: /sn:0 /dp:1 {0}(244,105)(348,105){1}
wire w4;    //: /sn:0 {0}(274,127)(293,127)(293,134)(303,134){1}
wire w2;    //: /sn:0 {0}(207,102)(215,102){1}
//: {2}(219,102)(223,102){3}
//: {4}(217,104)(217,129)(253,129){5}
wire w5;    //: /sn:0 {0}(273,150)(293,150)(293,139)(303,139){1}
//: enddecls

  //: joint g8 (Cin) @(213, 123) /w:[ 2 4 -1 1 ]
  //: output g4 (Cout) @(354,136) /sn:0 /w:[ 1 ]
  //: output g3 (S) @(345,105) /sn:0 /w:[ 1 ]
  //: input g2 (Cin) @(141,199) /sn:0 /w:[ 0 ]
  //: input g1 (B) @(141,173) /sn:0 /w:[ 0 ]
  and g10 (.I0(A), .I1(B), .Z(w5));   //: @(263,150) /sn:0 /tech:unit /w:[ 5 5 0 ]
  xor g6 (.I0(w2), .I1(Cin), .Z(S));   //: @(234,105) /sn:0 /delay:" 2" /w:[ 3 5 0 ]
  //: joint g9 (w2) @(217, 102) /w:[ 2 -1 1 4 ]
  and g7 (.I0(Cin), .I1(w2), .Z(w4));   //: @(264,127) /sn:0 /tech:unit /w:[ 3 5 0 ]
  //: joint g12 (B) @(161, 173) /w:[ 2 -1 1 4 ]
  //: joint g11 (A) @(152, 98) /w:[ 2 -1 1 4 ]
  xor g5 (.I0(A), .I1(B), .Z(w2));   //: @(197,102) /sn:0 /delay:" 2" /w:[ 3 3 0 ]
  //: input g0 (A) @(128,98) /sn:0 /w:[ 0 ]
  or g13 (.I0(w4), .I1(w5), .Z(Cout));   //: @(314,137) /sn:0 /tech:unit /w:[ 1 1 0 ]

endmodule
