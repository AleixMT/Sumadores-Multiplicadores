//: version "1.8.7"

module CarryLookahead_Logic(C3, P0, Cout, G0, P3, G1, P1, P2, C2, C1, G3, Cin, G2);
//: interface  /sz:(328, 96) /bd:[ Ti0>G0(286/328) Ti1>P0(267/328) Ti2>G1(210/328) Ti3>P1(189/328) Ti4>G2(139/328) Ti5>P2(117/328) Ti6>G3(55/328) Ti7>P3(28/328) Ri0>Cin(46/96) To0<C3(86/328) To1<C2(159/328) To2<C1(228/328) Lo0<Cout(39/96) ]
input G2;    //: /sn:0 {0}(49,313)(109,313)(109,301)(119,301){1}
input P1;    //: /sn:0 {0}(53,230)(109,230)(109,234)(119,234){1}
output C3;    //: /sn:0 /dp:1 {0}(360,293)(366,293)(366,292)(372,292){1}
//: {2}(376,292)(655,292)(655,289)(673,289){3}
//: {4}(374,294)(374,342)(391,342){5}
input G0;    //: /sn:0 {0}(74,187)(111,187)(111,169)(116,169){1}
output C2;    //: /sn:0 /dp:1 {0}(299,231)(320,231){1}
//: {2}(324,231)(610,231){3}
//: {4}(322,233)(322,290)(339,290){5}
input Cin;    //: /sn:0 {0}(85,65)(202,65)(202,162)(212,162){1}
input P3;    //: /sn:0 {0}(40,343)(112,343)(112,354)(122,354){1}
input G1;    //: /sn:0 {0}(51,249)(109,249)(109,239)(119,239){1}
output Cout;    //: /sn:0 /dp:1 {0}(412,345)(651,345)(651,376)(680,376){1}
input G3;    //: /sn:0 {0}(41,372)(112,372)(112,359)(122,359){1}
input P0;    //: /sn:0 {0}(75,145)(104,145)(104,164)(116,164){1}
output C1;    //: /sn:0 /dp:1 {0}(233,165)(263,165){1}
//: {2}(267,165)(609,165){3}
//: {4}(265,167)(265,228)(278,228){5}
input P2;    //: /sn:0 {0}(50,284)(109,284)(109,296)(119,296){1}
wire w6;    //: /sn:0 {0}(143,357)(382,357)(382,347)(391,347){1}
wire w4;    //: /sn:0 {0}(140,237)(268,237)(268,233)(278,233){1}
wire w3;    //: /sn:0 {0}(137,167)(212,167){1}
wire w5;    //: /sn:0 {0}(140,299)(329,299)(329,295)(339,295){1}
//: enddecls

  or g8 (.I0(P1), .I1(G1), .Z(w4));   //: @(130,237) /sn:0 /tech:unit /w:[ 1 1 0 ]
  and g4 (.I0(Cin), .I1(w3), .Z(C1));   //: @(223,165) /sn:0 /tech:unit /w:[ 1 1 0 ]
  and g16 (.I0(C2), .I1(w5), .Z(C3));   //: @(350,293) /sn:0 /tech:unit /w:[ 5 1 0 ]
  or g3 (.I0(P0), .I1(G0), .Z(w3));   //: @(127,167) /sn:0 /tech:unit /w:[ 1 1 0 ]
  //: output g17 (C3) @(670,289) /sn:0 /w:[ 3 ]
  //: input g2 (P0) @(73,145) /sn:0 /w:[ 0 ]
  //: output g23 (Cout) @(677,376) /sn:0 /w:[ 1 ]
  //: input g1 (G0) @(72,187) /sn:0 /w:[ 0 ]
  //: input g18 (P3) @(38,343) /sn:0 /w:[ 0 ]
  or g10 (.I0(P3), .I1(G3), .Z(w6));   //: @(133,357) /sn:0 /tech:unit /w:[ 1 1 0 ]
  //: input g6 (G1) @(49,249) /sn:0 /w:[ 0 ]
  or g9 (.I0(P2), .I1(G2), .Z(w5));   //: @(130,299) /sn:0 /tech:unit /w:[ 1 1 0 ]
  //: input g7 (P1) @(51,230) /sn:0 /w:[ 0 ]
  //: joint g22 (C3) @(374, 292) /w:[ 2 -1 1 4 ]
  //: input g12 (P2) @(48,284) /sn:0 /w:[ 0 ]
  and g14 (.I0(C1), .I1(w4), .Z(C2));   //: @(289,231) /sn:0 /tech:unit /w:[ 5 1 0 ]
  //: output g11 (C2) @(607,231) /sn:0 /w:[ 3 ]
  //: output g5 (C1) @(606,165) /sn:0 /w:[ 3 ]
  and g21 (.I0(C3), .I1(w6), .Z(Cout));   //: @(402,345) /sn:0 /tech:unit /w:[ 5 1 0 ]
  //: input g19 (G3) @(39,372) /sn:0 /w:[ 0 ]
  //: joint g20 (C2) @(322, 231) /w:[ 2 -1 1 4 ]
  //: joint g15 (C1) @(265, 165) /w:[ 2 -1 1 4 ]
  //: input g0 (Cin) @(83,65) /sn:0 /w:[ 0 ]
  //: input g13 (G2) @(47,313) /sn:0 /w:[ 0 ]

endmodule

module PFA_v1(C, B, P, S, A, G);
//: interface  /sz:(126, 115) /bd:[ Ti0>A(21/126) Ti1>B(82/126) Ri0>C(56/115) Bo0<S(99/126) Bo1<P(11/126) Bo2<G(56/126) ]
input B;    //: /sn:0 {0}(144,200)(161,200){1}
//: {2}(165,200)(202,200)(202,177)(210,177){3}
//: {4}(163,202)(163,320){5}
//: {6}(165,322)(231,322){7}
//: {8}(163,324)(163,361)(240,361){9}
input A;    //: /sn:0 {0}(151,147)(178,147){1}
//: {2}(182,147)(202,147)(202,172)(210,172){3}
//: {4}(180,149)(180,317)(188,317){5}
//: {6}(192,317)(231,317){7}
//: {8}(190,319)(190,356)(240,356){9}
output G;    //: /sn:0 /dp:1 {0}(261,359)(337,359)(337,385)(346,385){1}
input C;    //: /sn:0 {0}(149,271)(266,271)(266,186)(276,186){1}
output P;    //: /sn:0 /dp:1 {0}(252,320)(312,320)(312,319)(322,319){1}
output S;    //: /sn:0 /dp:1 {0}(297,184)(394,184)(394,198)(406,198){1}
wire w2;    //: /sn:0 {0}(231,175)(267,175)(267,181)(276,181){1}
//: enddecls

  xor g4 (.I0(w2), .I1(C), .Z(S));   //: @(287,184) /sn:0 /delay:" 2" /w:[ 1 1 0 ]
  //: joint g8 (B) @(163, 200) /w:[ 2 -1 1 4 ]
  xor g3 (.I0(A), .I1(B), .Z(w2));   //: @(221,175) /sn:0 /delay:" 2" /w:[ 3 3 0 ]
  //: input g2 (C) @(147,271) /sn:0 /w:[ 0 ]
  //: input g1 (B) @(142,200) /sn:0 /w:[ 0 ]
  and g10 (.I0(A), .I1(B), .Z(G));   //: @(251,359) /sn:0 /delay:" 1" /w:[ 9 9 0 ]
  or g6 (.I0(A), .I1(B), .Z(P));   //: @(242,320) /sn:0 /delay:" 1" /w:[ 7 7 0 ]
  //: joint g7 (A) @(180, 147) /w:[ 2 -1 1 4 ]
  //: output g9 (P) @(319,319) /sn:0 /w:[ 1 ]
  //: joint g12 (A) @(190, 317) /w:[ 6 -1 5 8 ]
  //: output g5 (S) @(403,198) /sn:0 /w:[ 1 ]
  //: joint g11 (B) @(163, 322) /w:[ 6 5 -1 8 ]
  //: input g0 (A) @(149,147) /sn:0 /w:[ 0 ]
  //: output g13 (G) @(343,385) /sn:0 /w:[ 1 ]

endmodule

module main;    //: root_module
wire w13;    //: /sn:0 {0}(-480,528)(-480,576){1}
//: {2}(-478,578)(-462,578)(-462,565){3}
//: {4}(-480,580)(-480,611)(-492,611)(-492,651){5}
wire w6;    //: /sn:0 {0}(-279,526)(-279,578)(-338,578)(-338,597){1}
//: {2}(-336,599)(-313,599)(-313,611)(-298,611)(-298,601){3}
//: {4}(-338,601)(-338,638)(-340,638)(-340,651){5}
wire w16;    //: /sn:0 {0}(196,256)(196,322){1}
//: {2}(198,324)(228,324)(228,322){3}
//: {4}(196,326)(196,371)(217,371)(217,379){5}
wire w7;    //: /sn:0 {0}(-1943,949)(-1943,982)(-1945,982)(-1945,1015){1}
//: {2}(-1943,1017)(-1877,1017)(-1877,1051)(-1861,1051)(-1861,1041){3}
//: {4}(-1945,1019)(-1945,1066)(-2005,1066)(-2005,1074){5}
wire w65;    //: /sn:0 {0}(-1483,602)(-1478,602)(-1478,628){1}
wire w58;    //: /sn:0 {0}(-1661,736)(-1661,782){1}
//: {2}(-1659,784)(-1635,784)(-1635,777){3}
//: {4}(-1661,786)(-1661,860)(-1640,860)(-1640,868){5}
wire w88;    //: /sn:0 {0}(-2441,942)(-2441,990)(-2425,990)(-2425,980){1}
wire w50;    //: /sn:0 {0}(-1666,588)(-1651,588)(-1651,619){1}
wire w34;    //: /sn:0 {0}(299,379)(299,351)(332,351)(332,196)(326,196){1}
//: {2}(324,194)(324,184)(323,184)(323,173){3}
//: {4}(322,196)(312,196){5}
wire w81;    //: /sn:0 {0}(-2529,942)(-2529,988){1}
//: {2}(-2527,990)(-2503,990)(-2503,983){3}
//: {4}(-2529,992)(-2529,1066)(-2508,1066)(-2508,1074){5}
wire w59;    //: /sn:0 {0}(-1054,915)(-958,915)(-958,683)(-960,683){1}
//: {2}(-962,681)(-962,678)(-894,678){3}
//: {4}(-892,676)(-892,657){5}
//: {6}(-892,680)(-892,691)(-861,691){7}
//: {8}(-964,683)(-1004,683){9}
wire w72;    //: /sn:0 {0}(-1120,609)(-1110,609)(-1110,626){1}
wire w62;    //: /sn:0 {0}(-1250,868)(-1250,833)(-1180,833)(-1180,687){1}
//: {2}(-1180,683)(-1180,673)(-1186,673)(-1186,643){3}
//: {4}(-1182,685)(-1198,685){5}
wire w39;    //: /sn:0 {0}(-416,651)(-416,616)(-346,616)(-346,470){1}
//: {2}(-346,466)(-346,456)(-352,456)(-352,426){3}
//: {4}(-348,468)(-364,468){5}
wire w4;    //: /sn:0 {0}(571,254)(571,306)(512,306)(512,325){1}
//: {2}(514,327)(537,327)(537,339)(552,339)(552,329){3}
//: {4}(512,329)(512,366)(510,366)(510,379){5}
wire w25;    //: /sn:0 {0}(564,120)(574,120)(574,137){1}
wire w56;    //: /sn:0 {0}(-1488,745)(-1488,811){1}
//: {2}(-1486,813)(-1456,813)(-1456,811){3}
//: {4}(-1488,815)(-1488,860)(-1467,860)(-1467,868){5}
wire w82;    //: /sn:0 {0}(-1922,1121)(-1826,1121)(-1826,891){1}
//: {2}(-1824,889)(-1738,889)(-1738,890)(-1728,890){3}
//: {4}(-1726,888)(-1726,874){5}
//: {6}(-1726,892)(-1726,908)(-1695,908){7}
//: {8}(-1828,889)(-1872,889){9}
wire w36;    //: /sn:0 {0}(-220,698)(-121,698)(-121,468){1}
//: {2}(-119,466)(-54,466)(-54,412)(-44,412){3}
//: {4}(-42,410)(-42,385){5}
//: {6}(-42,414)(-42,419)(-11,419){7}
//: {8}(-123,466)(-170,466){9}
wire w3;    //: /sn:0 {0}(609,254)(609,287)(607,287)(607,320){1}
//: {2}(609,322)(675,322)(675,356)(691,356)(691,346){3}
//: {4}(607,324)(607,371)(547,371)(547,379){5}
wire w22;    //: /sn:0 {0}(23,247)(23,293){1}
//: {2}(25,295)(49,295)(49,288){3}
//: {4}(23,297)(23,371)(44,371)(44,379){5}
wire w0;    //: /sn:0 /dp:1 {0}(439,289)(439,299)(458,299)(458,256){1}
wire w60;    //: /sn:0 {0}(-1527,868)(-1527,689)(-1528,689)(-1528,678){1}
//: {2}(-1528,674)(-1528,664)(-1534,664)(-1534,631){3}
//: {4}(-1530,676)(-1545,676){5}
wire w20;    //: /sn:0 {0}(377,112)(380,112)(380,139){1}
wire w71;    //: /sn:0 {0}(-1045,784)(-1045,794)(-1032,794)(-1032,743){1}
wire w30;    //: /sn:0 {0}(-827,519)(-827,565){1}
//: {2}(-825,567)(-801,567)(-801,560){3}
//: {4}(-827,569)(-827,643)(-806,643)(-806,651){5}
wire w29;    //: /sn:0 {0}(-782,519)(-782,598){1}
//: {2}(-780,600)(-746,600)(-746,586){3}
//: {4}(-782,602)(-782,643)(-753,643)(-753,651){5}
wire w42;    //: /sn:0 {0}(-593,390)(-583,390)(-583,411){1}
wire w37;    //: /sn:0 {0}(-693,651)(-693,472)(-694,472)(-694,461){1}
//: {2}(-694,457)(-694,447)(-700,447)(-700,414){3}
//: {4}(-696,459)(-711,459){5}
wire w73;    //: /sn:0 {0}(-1063,602)(-1049,602)(-1049,626){1}
wire w66;    //: /sn:0 {0}(-1427,607)(-1417,607)(-1417,628){1}
wire w12;    //: /sn:0 {0}(-435,528)(-435,571)(-449,571)(-449,606){1}
//: {2}(-447,608)(-441,608)(-441,621)(-426,621)(-426,611){3}
//: {4}(-449,610)(-449,642)(-451,642)(-451,651){5}
wire w18;    //: /sn:0 {0}(201,113)(206,113)(206,139){1}
wire w19;    //: /sn:0 {0}(257,118)(267,118)(267,139){1}
wire w63;    //: /sn:0 {0}(-1599,588)(-1590,588)(-1590,619){1}
wire w10;    //: /sn:0 {0}(370,256)(370,304){1}
//: {2}(372,306)(388,306)(388,293){3}
//: {4}(370,308)(370,339)(358,339)(358,379){5}
wire w23;    //: /sn:0 {0}(111,247)(111,295)(127,295)(127,285){1}
wire w91;    //: /sn:0 {0}(-2268,951)(-2268,995)(-2248,995)(-2248,985){1}
wire w84;    //: /sn:0 {0}(-2253,1074)(-2253,1046)(-2220,1046)(-2220,891)(-2226,891){1}
//: {2}(-2228,889)(-2228,879)(-2229,879)(-2229,868){3}
//: {4}(-2230,891)(-2240,891){5}
wire w70;    //: /sn:0 {0}(-1256,595)(-1243,595)(-1243,628){1}
wire w54;    //: /sn:0 {0}(-1314,745)(-1314,793){1}
//: {2}(-1312,795)(-1296,795)(-1296,782){3}
//: {4}(-1314,797)(-1314,828)(-1326,828)(-1326,868){5}
wire w86;    //: /sn:0 {0}(-2594,1080)(-2594,1114)(-2563,1114){1}
wire w21;    //: /sn:0 {0}(68,247)(68,326){1}
//: {2}(70,328)(104,328)(104,314){3}
//: {4}(68,330)(68,371)(97,371)(97,379){5}
wire w24;    //: /sn:0 {0}(428,106)(441,106)(441,139){1}
wire w31;    //: /sn:0 {0}(-765,371)(-756,371)(-756,402){1}
wire w1;    //: /sn:0 /dp:1 {0}(639,295)(639,305)(652,305)(652,254){1}
wire w68;    //: /sn:0 {0}(-1245,778)(-1245,788)(-1226,788)(-1226,745){1}
wire w32;    //: /sn:0 {0}(630,426)(726,426)(726,194){1}
//: {2}(726,190)(726,163)(715,163){3}
//: {4}(724,192)(688,192)(688,194)(680,194){5}
wire w53;    //: /sn:0 {0}(-1269,745)(-1269,788)(-1283,788)(-1283,823){1}
//: {2}(-1281,825)(-1275,825)(-1275,838)(-1260,838)(-1260,828){3}
//: {4}(-1283,827)(-1283,859)(-1285,859)(-1285,868){5}
wire w46;    //: /sn:0 {0}(-422,378)(-409,378)(-409,411){1}
wire w8;    //: /sn:0 {0}(18,99)(33,99)(33,130){1}
wire w95;    //: /sn:0 {0}(-1913,990)(-1913,1000)(-1900,1000)(-1900,949){1}
wire w89;    //: /sn:0 {0}(-2351,808)(-2346,808)(-2346,834){1}
wire w52;    //: /sn:0 {0}(-1113,743)(-1113,795)(-1172,795)(-1172,814){1}
//: {2}(-1170,816)(-1147,816)(-1147,828)(-1132,828)(-1132,818){3}
//: {4}(-1172,818)(-1172,855)(-1174,855)(-1174,868){5}
wire w75;    //: /sn:0 {0}(-1981,949)(-1981,1001)(-2040,1001)(-2040,1020){1}
//: {2}(-2038,1022)(-2015,1022)(-2015,1034)(-2000,1034)(-2000,1024){3}
//: {4}(-2040,1024)(-2040,1061)(-2042,1061)(-2042,1074){5}
wire w44;    //: /sn:0 {0}(-411,561)(-411,571)(-392,571)(-392,528){1}
wire w27;    //: /sn:0 {0}(-609,528)(-609,569){1}
//: {2}(-607,571)(-593,571)(-593,578)(-578,578)(-578,568){3}
//: {4}(-609,573)(-609,625)(-590,625)(-590,651){5}
wire w17;    //: /sn:0 {0}(284,256)(284,300)(304,300)(304,290){1}
wire w80;    //: /sn:0 {0}(-2484,942)(-2484,1021){1}
//: {2}(-2482,1023)(-2448,1023)(-2448,1009){3}
//: {4}(-2484,1025)(-2484,1066)(-2455,1066)(-2455,1074){5}
wire w67;    //: /sn:0 {0}(-1400,745)(-1400,789)(-1380,789)(-1380,779){1}
wire w28;    //: /sn:0 {0}(-654,528)(-654,594){1}
//: {2}(-652,596)(-622,596)(-622,594){3}
//: {4}(-654,598)(-654,643)(-633,643)(-633,651){5}
wire w33;    //: /sn:0 {0}(434,379)(434,344)(504,344)(504,198){1}
//: {2}(504,194)(504,184)(498,184)(498,154){3}
//: {4}(502,196)(486,196){5}
wire w35;    //: /sn:0 {0}(157,379)(157,200)(156,200)(156,189){1}
//: {2}(156,185)(156,175)(150,175)(150,142){3}
//: {4}(154,187)(139,187){5}
wire w69;    //: /sn:0 {0}(-1307,601)(-1304,601)(-1304,628){1}
wire w49;    //: /sn:0 {0}(-229,385)(-215,385)(-215,409){1}
wire w45;    //: /sn:0 {0}(-473,384)(-470,384)(-470,411){1}
wire w14;    //: /sn:0 {0}(85,99)(94,99)(94,130){1}
wire w78;    //: /sn:0 {0}(-2311,951)(-2311,992){1}
//: {2}(-2309,994)(-2295,994)(-2295,1001)(-2280,1001)(-2280,991){3}
//: {4}(-2311,996)(-2311,1048)(-2292,1048)(-2292,1074){5}
wire w74;    //: /sn:0 {0}(-2534,794)(-2519,794)(-2519,825){1}
wire w48;    //: /sn:0 {0}(-286,392)(-276,392)(-276,409){1}
wire w41;    //: /sn:0 {0}(-649,385)(-644,385)(-644,411){1}
wire w11;    //: /sn:0 {0}(-832,371)(-817,371)(-817,402){1}
wire w47;    //: /sn:0 {0}(-211,567)(-211,577)(-198,577)(-198,526){1}
wire w90;    //: /sn:0 {0}(-2295,813)(-2285,813)(-2285,834){1}
wire w85;    //: /sn:0 {0}(-2118,1074)(-2118,1039)(-2048,1039)(-2048,893){1}
//: {2}(-2048,889)(-2048,879)(-2054,879)(-2054,849){3}
//: {4}(-2050,891)(-2066,891){5}
wire w83;    //: /sn:0 {0}(-2395,1074)(-2395,895)(-2396,895)(-2396,884){1}
//: {2}(-2396,880)(-2396,870)(-2402,870)(-2402,837){3}
//: {4}(-2398,882)(-2413,882){5}
wire w15;    //: /sn:0 {0}(241,256)(241,297){1}
//: {2}(243,299)(257,299)(257,306)(272,306)(272,296){3}
//: {4}(241,301)(241,353)(260,353)(260,379){5}
wire w94;    //: /sn:0 {0}(-2124,801)(-2111,801)(-2111,834){1}
wire w92;    //: /sn:0 {0}(-2113,984)(-2113,994)(-2094,994)(-2094,951){1}
wire w61;    //: /sn:0 {0}(-1385,868)(-1385,840)(-1352,840)(-1352,685)(-1358,685){1}
//: {2}(-1360,683)(-1360,673)(-1361,673)(-1361,662){3}
//: {4}(-1362,685)(-1372,685){5}
wire w55;    //: /sn:0 {0}(-1443,745)(-1443,786){1}
//: {2}(-1441,788)(-1427,788)(-1427,795)(-1412,795)(-1412,785){3}
//: {4}(-1443,790)(-1443,842)(-1424,842)(-1424,868){5}
wire w38;    //: /sn:0 {0}(-551,651)(-551,623)(-518,623)(-518,468)(-524,468){1}
//: {2}(-526,466)(-526,456)(-527,456)(-527,445){3}
//: {4}(-528,468)(-538,468){5}
wire w5;    //: /sn:0 {0}(-241,526)(-241,559)(-243,559)(-243,592){1}
//: {2}(-241,594)(-175,594)(-175,628)(-159,628)(-159,618){3}
//: {4}(-243,596)(-243,643)(-303,643)(-303,651){5}
wire w87;    //: /sn:0 {0}(-2467,794)(-2458,794)(-2458,825){1}
wire w64;    //: /sn:0 {0}(-1573,736)(-1573,784)(-1557,784)(-1557,774){1}
wire w43;    //: /sn:0 {0}(-566,528)(-566,572)(-546,572)(-546,562){1}
wire w97;    //: /sn:0 {0}(-1931,808)(-1917,808)(-1917,832){1}
wire w96;    //: /sn:0 {0}(-1988,815)(-1978,815)(-1978,832){1}
wire w76;    //: /sn:0 {0}(-2137,951)(-2137,994)(-2151,994)(-2151,1029){1}
//: {2}(-2149,1031)(-2143,1031)(-2143,1044)(-2128,1044)(-2128,1034){3}
//: {4}(-2151,1033)(-2151,1065)(-2153,1065)(-2153,1074){5}
wire w9;    //: /sn:0 {0}(415,256)(415,299)(401,299)(401,334){1}
//: {2}(403,336)(409,336)(409,349)(424,349)(424,339){3}
//: {4}(401,338)(401,370)(399,370)(399,379){5}
wire w26;    //: /sn:0 {0}(621,113)(635,113)(635,137){1}
wire w93;    //: /sn:0 {0}(-2175,807)(-2172,807)(-2172,834){1}
wire w79;    //: /sn:0 {0}(-2356,951)(-2356,1017){1}
//: {2}(-2354,1019)(-2324,1019)(-2324,1017){3}
//: {4}(-2356,1021)(-2356,1066)(-2335,1066)(-2335,1074){5}
wire w77;    //: /sn:0 {0}(-2182,951)(-2182,999){1}
//: {2}(-2180,1001)(-2164,1001)(-2164,988){3}
//: {4}(-2182,1003)(-2182,1034)(-2194,1034)(-2194,1074){5}
wire w57;    //: /sn:0 {0}(-1616,736)(-1616,815){1}
//: {2}(-1614,817)(-1580,817)(-1580,803){3}
//: {4}(-1616,819)(-1616,860)(-1587,860)(-1587,868){5}
wire w51;    //: /sn:0 {0}(-1075,743)(-1075,776)(-1077,776)(-1077,809){1}
//: {2}(-1075,811)(-1009,811)(-1009,845)(-993,845)(-993,835){3}
//: {4}(-1077,813)(-1077,860)(-1137,860)(-1137,868){5}
wire w40;    //: /sn:0 {0}(-739,519)(-739,567)(-723,567)(-723,557){1}
//: enddecls

  PFA_v1 g164 (.A(w96), .B(w97), .C(w82), .S(w95), .P(w75), .G(w7));   //: @(-1999, 833) /sz:(126, 115) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>9 Bo0<1 Bo1<0 Bo2<0 ]
  //: switch g8 (w8) @(1,99) /sn:0 /w:[ 0 ] /st:1
  CarryLookahead_Logic g4 (.G0(w3), .P0(w4), .G1(w9), .P1(w10), .G2(w15), .P2(w16), .G3(w21), .P3(w22), .Cin(w32), .C3(w35), .C2(w34), .C1(w33), .Cout(w36));   //: @(-10, 380) /sz:(639, 96) /sn:0 /p:[ Ti0>5 Ti1>5 Ti2>5 Ti3>5 Ti4>5 Ti5>5 Ti6>5 Ti7>5 Ri0>0 To0<0 To1<0 To2<0 Lo0<7 ]
  //: joint g116 (w60) @(-1528, 676) /w:[ -1 2 4 1 ]
  //: joint g157 (w82) @(-1726, 890) /w:[ -1 4 3 6 ]
  //: joint g17 (w33) @(504, 196) /w:[ -1 2 4 1 ]
  PFA_v1 g137 (.A(w93), .B(w94), .C(w85), .S(w92), .P(w77), .G(w76));   //: @(-2193, 835) /sz:(126, 115) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>5 Bo0<1 Bo1<0 Bo2<0 ]
  led g30 (.I(w9));   //: @(424,332) /sn:0 /w:[ 3 ] /type:0
  //: joint g74 (w37) @(-694, 459) /w:[ -1 2 4 1 ]
  led g92 (.I(w53));   //: @(-1260,821) /sn:0 /w:[ 3 ] /type:0
  PFA_v1 g130 (.A(w74), .B(w87), .C(w83), .S(w88), .P(w81), .G(w80));   //: @(-2540, 826) /sz:(126, 115) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>5 Bo0<0 Bo1<0 Bo2<0 ]
  PFA_v1 g1 (.A(w20), .B(w24), .C(w33), .S(w0), .P(w10), .G(w9));   //: @(359, 140) /sz:(126, 115) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>5 Bo0<1 Bo1<0 Bo2<0 ]
  led g77 (.I(w13));   //: @(-462,558) /sn:0 /w:[ 3 ] /type:0
  led g111 (.I(w52));   //: @(-1132,811) /sn:0 /w:[ 3 ] /type:0
  led g144 (.I(w86));   //: @(-2594,1073) /sn:0 /w:[ 0 ] /type:0
  led g51 (.I(w44));   //: @(-411,554) /sn:0 /w:[ 0 ] /type:0
  led g161 (.I(w77));   //: @(-2164,981) /sn:0 /w:[ 3 ] /type:0
  led g70 (.I(w27));   //: @(-578,561) /sn:0 /w:[ 3 ] /type:0
  led g149 (.I(w79));   //: @(-2324,1010) /sn:0 /w:[ 3 ] /type:0
  led g25 (.I(w1));   //: @(639,288) /sn:0 /w:[ 0 ] /type:0
  //: switch g10 (w18) @(184,113) /sn:0 /w:[ 0 ] /st:1
  led g65 (.I(w28));   //: @(-622,587) /sn:0 /w:[ 3 ] /type:0
  //: joint g103 (w55) @(-1443, 788) /w:[ 2 1 -1 4 ]
  //: joint g64 (w13) @(-480, 578) /w:[ 2 1 -1 4 ]
  PFA_v1 g49 (.A(w41), .B(w42), .C(w38), .S(w43), .P(w28), .G(w27));   //: @(-665, 412) /sz:(126, 115) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>5 Bo0<0 Bo1<0 Bo2<0 ]
  //: switch g72 (w42) @(-610,390) /sn:0 /w:[ 0 ] /st:0
  //: joint g142 (w82) @(-1826, 889) /w:[ 2 -1 8 1 ]
  //: joint g136 (w80) @(-2484, 1023) /w:[ 2 1 -1 4 ]
  //: joint g6 (w32) @(726, 192) /w:[ -1 2 4 1 ]
  led g7 (.I(w36));   //: @(-42,378) /sn:0 /w:[ 5 ] /type:0
  //: joint g35 (w15) @(241, 299) /w:[ 2 1 -1 4 ]
  led g56 (.I(w47));   //: @(-211,560) /sn:0 /w:[ 0 ] /type:0
  //: joint g58 (w36) @(-121, 466) /w:[ 2 -1 8 1 ]
  //: joint g124 (w56) @(-1488, 813) /w:[ 2 1 -1 4 ]
  led g98 (.I(w71));   //: @(-1045,777) /sn:0 /w:[ 0 ] /type:0
  led g67 (.I(w30));   //: @(-801,553) /sn:0 /w:[ 3 ] /type:0
  led g85 (.I(w62));   //: @(-1186,636) /sn:0 /w:[ 3 ] /type:0
  //: switch g126 (w74) @(-2551,794) /sn:0 /w:[ 0 ] /st:1
  //: joint g33 (w10) @(370, 306) /w:[ 2 1 -1 4 ]
  //: joint g54 (w6) @(-338, 599) /w:[ 2 1 -1 4 ]
  led g40 (.I(w22));   //: @(49,281) /sn:0 /w:[ 3 ] /type:0
  //: joint g52 (w29) @(-782, 600) /w:[ 2 1 -1 4 ]
  //: joint g81 (w5) @(-243, 594) /w:[ 2 1 -1 4 ]
  led g163 (.I(w80));   //: @(-2448,1002) /sn:0 /w:[ 3 ] /type:0
  led g132 (.I(w91));   //: @(-2248,978) /sn:0 /w:[ 1 ] /type:0
  //: switch g12 (w20) @(360,112) /sn:0 /w:[ 0 ] /st:0
  //: joint g108 (w58) @(-1661, 784) /w:[ 2 1 -1 4 ]
  led g131 (.I(w7));   //: @(-1861,1034) /sn:0 /w:[ 3 ] /type:0
  //: joint g106 (w54) @(-1314, 795) /w:[ 2 1 -1 4 ]
  //: joint g96 (w52) @(-1172, 816) /w:[ 2 1 -1 4 ]
  //: joint g19 (w34) @(324, 196) /w:[ 1 2 4 -1 ]
  //: switch g114 (w66) @(-1444,607) /sn:0 /w:[ 0 ] /st:0
  //: joint g117 (w61) @(-1360, 685) /w:[ 1 2 4 -1 ]
  //: switch g78 (w49) @(-246,385) /sn:0 /w:[ 0 ] /st:1
  //: switch g125 (w70) @(-1273,595) /sn:0 /w:[ 0 ] /st:1
  //: switch g155 (w96) @(-2005,815) /sn:0 /w:[ 0 ] /st:0
  //: joint g63 (w12) @(-449, 608) /w:[ 2 1 -1 4 ]
  led g93 (.I(w68));   //: @(-1245,771) /sn:0 /w:[ 0 ] /type:0
  //: joint g105 (w53) @(-1283, 825) /w:[ 2 1 -1 4 ]
  //: switch g113 (w72) @(-1137,609) /sn:0 /w:[ 0 ] /st:0
  //: joint g100 (w59) @(-962, 683) /w:[ 1 2 8 -1 ]
  PFA_v1 g0 (.A(w25), .B(w26), .C(w32), .S(w1), .P(w4), .G(w3));   //: @(553, 138) /sz:(126, 115) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>5 Bo0<1 Bo1<0 Bo2<0 ]
  led g38 (.I(w21));   //: @(104,307) /sn:0 /w:[ 3 ] /type:0
  led g43 (.I(w39));   //: @(-352,419) /sn:0 /w:[ 3 ] /type:0
  //: switch g101 (w63) @(-1616,588) /sn:0 /w:[ 0 ] /st:1
  led g48 (.I(w43));   //: @(-546,555) /sn:0 /w:[ 1 ] /type:0
  //: joint g37 (w16) @(196, 324) /w:[ 2 1 -1 4 ]
  PFA_v1 g80 (.A(w48), .B(w49), .C(w36), .S(w47), .P(w6), .G(w5));   //: @(-297, 410) /sz:(126, 115) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>9 Bo0<1 Bo1<0 Bo2<0 ]
  PFA_v1 g95 (.A(w69), .B(w70), .C(w62), .S(w68), .P(w54), .G(w53));   //: @(-1325, 629) /sz:(126, 115) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>5 Bo0<1 Bo1<0 Bo2<0 ]
  //: switch g120 (w73) @(-1080,602) /sn:0 /w:[ 0 ] /st:1
  PFA_v1 g122 (.A(w72), .B(w73), .C(w59), .S(w71), .P(w52), .G(w51));   //: @(-1131, 627) /sz:(126, 115) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>9 Bo0<1 Bo1<0 Bo2<0 ]
  led g76 (.I(w37));   //: @(-700,407) /sn:0 /w:[ 3 ] /type:0
  //: switch g152 (w93) @(-2192,807) /sn:0 /w:[ 0 ] /st:0
  CarryLookahead_Logic g44 (.G0(w5), .P0(w6), .G1(w12), .P1(w13), .G2(w27), .P2(w28), .G3(w29), .P3(w30), .Cin(w36), .C3(w37), .C2(w38), .C1(w39), .Cout(w59));   //: @(-860, 652) /sz:(639, 96) /sn:0 /p:[ Ti0>5 Ti1>5 Ti2>5 Ti3>5 Ti4>5 Ti5>5 Ti6>5 Ti7>5 Ri0>0 To0<0 To1<0 To2<0 Lo0<7 ]
  //: joint g75 (w38) @(-526, 468) /w:[ 1 2 4 -1 ]
  //: joint g159 (w84) @(-2228, 891) /w:[ 1 2 4 -1 ]
  led g16 (.I(w33));   //: @(498,147) /sn:0 /w:[ 3 ] /type:0
  PFA_v1 g3 (.A(w8), .B(w14), .C(w35), .S(w23), .P(w22), .G(w21));   //: @(12, 131) /sz:(126, 115) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>5 Bo0<0 Bo1<0 Bo2<0 ]
  led g47 (.I(w5));   //: @(-159,611) /sn:0 /w:[ 3 ] /type:0
  //: switch g143 (w87) @(-2484,794) /sn:0 /w:[ 0 ] /st:1
  led g26 (.I(w3));   //: @(691,339) /sn:0 /w:[ 3 ] /type:0
  led g90 (.I(w67));   //: @(-1380,772) /sn:0 /w:[ 1 ] /type:0
  led g109 (.I(w58));   //: @(-1635,770) /sn:0 /w:[ 3 ] /type:0
  //: joint g158 (w83) @(-2396, 882) /w:[ -1 2 4 1 ]
  PFA_v1 g2 (.A(w18), .B(w19), .C(w34), .S(w17), .P(w16), .G(w15));   //: @(185, 140) /sz:(126, 115) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>5 Bo0<0 Bo1<0 Bo2<0 ]
  CarryLookahead_Logic g128 (.G0(w7), .P0(w75), .G1(w76), .P1(w77), .G2(w78), .P2(w79), .G3(w80), .P3(w81), .Cin(w82), .C3(w83), .C2(w84), .C1(w85), .Cout(w86));   //: @(-2562, 1075) /sz:(639, 96) /sn:0 /p:[ Ti0>5 Ti1>5 Ti2>5 Ti3>5 Ti4>5 Ti5>5 Ti6>5 Ti7>5 Ri0>0 To0<0 To1<0 To2<0 Lo0<1 ]
  led g23 (.I(w17));   //: @(304,283) /sn:0 /w:[ 1 ] /type:0
  PFA_v1 g91 (.A(w65), .B(w66), .C(w61), .S(w67), .P(w56), .G(w55));   //: @(-1499, 629) /sz:(126, 115) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>5 Bo0<0 Bo1<0 Bo2<0 ]
  //: switch g141 (w89) @(-2368,808) /sn:0 /w:[ 0 ] /st:1
  led g24 (.I(w0));   //: @(439,282) /sn:0 /w:[ 0 ] /type:0
  //: joint g39 (w21) @(68, 328) /w:[ 2 1 -1 4 ]
  CarryLookahead_Logic g86 (.G0(w51), .P0(w52), .G1(w53), .P1(w54), .G2(w55), .P2(w56), .G3(w57), .P3(w58), .Cin(w59), .C3(w60), .C2(w61), .C1(w62), .Cout(w82));   //: @(-1694, 869) /sz:(639, 96) /sn:0 /p:[ Ti0>5 Ti1>5 Ti2>5 Ti3>5 Ti4>5 Ti5>5 Ti6>5 Ti7>5 Ri0>0 To0<0 To1<0 To2<0 Lo0<7 ]
  led g104 (.I(w64));   //: @(-1557,767) /sn:0 /w:[ 1 ] /type:0
  led g127 (.I(w85));   //: @(-2054,842) /sn:0 /w:[ 3 ] /type:0
  //: joint g29 (w4) @(512, 327) /w:[ 2 1 -1 4 ]
  led g60 (.I(w59));   //: @(-892,650) /sn:0 /w:[ 5 ] /type:0
  //: switch g110 (w69) @(-1324,601) /sn:0 /w:[ 0 ] /st:0
  led g121 (.I(w57));   //: @(-1580,796) /sn:0 /w:[ 3 ] /type:0
  led g18 (.I(w34));   //: @(323,166) /sn:0 /w:[ 3 ] /type:0
  //: joint g82 (w28) @(-654, 596) /w:[ 2 1 -1 4 ]
  //: joint g94 (w57) @(-1616, 817) /w:[ 2 1 -1 4 ]
  led g119 (.I(w54));   //: @(-1296,775) /sn:0 /w:[ 3 ] /type:0
  //: joint g166 (w79) @(-2356, 1019) /w:[ 2 1 -1 4 ]
  led g154 (.I(w78));   //: @(-2280,984) /sn:0 /w:[ 3 ] /type:0
  led g107 (.I(w56));   //: @(-1456,804) /sn:0 /w:[ 3 ] /type:0
  led g50 (.I(w12));   //: @(-426,604) /sn:0 /w:[ 3 ] /type:0
  PFA_v1 g133 (.A(w89), .B(w90), .C(w84), .S(w91), .P(w79), .G(w78));   //: @(-2367, 835) /sz:(126, 115) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>5 Bo0<0 Bo1<0 Bo2<0 ]
  //: switch g9 (w14) @(68,99) /sn:0 /w:[ 0 ] /st:1
  //: switch g68 (w45) @(-490,384) /sn:0 /w:[ 0 ] /st:0
  //: joint g73 (w36) @(-42, 412) /w:[ -1 4 3 6 ]
  led g22 (.I(w23));   //: @(127,278) /sn:0 /w:[ 1 ] /type:0
  //: joint g31 (w9) @(401, 336) /w:[ 2 1 -1 4 ]
  //: switch g59 (w31) @(-782,371) /sn:0 /w:[ 0 ] /st:1
  //: switch g71 (w48) @(-303,392) /sn:0 /w:[ 0 ] /st:0
  led g102 (.I(w82));   //: @(-1726,867) /sn:0 /w:[ 5 ] /type:0
  //: joint g87 (w62) @(-1180, 685) /w:[ -1 2 4 1 ]
  //: switch g83 (w46) @(-439,378) /sn:0 /w:[ 0 ] /st:1
  //: switch g99 (w65) @(-1500,602) /sn:0 /w:[ 0 ] /st:1
  led g36 (.I(w16));   //: @(228,315) /sn:0 /w:[ 3 ] /type:0
  //: joint g41 (w22) @(23, 295) /w:[ 2 1 -1 4 ]
  //: joint g45 (w39) @(-346, 468) /w:[ -1 2 4 1 ]
  //: switch g156 (w90) @(-2312,813) /sn:0 /w:[ 0 ] /st:0
  //: joint g138 (w75) @(-2040, 1022) /w:[ 2 1 -1 4 ]
  //: switch g42 (w11) @(-849,371) /sn:0 /w:[ 0 ] /st:1
  led g69 (.I(w6));   //: @(-298,594) /sn:0 /w:[ 3 ] /type:0
  //: switch g167 (w94) @(-2141,801) /sn:0 /w:[ 0 ] /st:1
  led g151 (.I(w81));   //: @(-2503,976) /sn:0 /w:[ 3 ] /type:0
  //: joint g66 (w30) @(-827, 567) /w:[ 2 1 -1 4 ]
  //: switch g162 (w97) @(-1948,808) /sn:0 /w:[ 0 ] /st:1
  led g153 (.I(w75));   //: @(-2000,1017) /sn:0 /w:[ 3 ] /type:0
  led g146 (.I(w88));   //: @(-2425,973) /sn:0 /w:[ 1 ] /type:0
  led g28 (.I(w4));   //: @(552,322) /sn:0 /w:[ 3 ] /type:0
  led g34 (.I(w15));   //: @(272,289) /sn:0 /w:[ 3 ] /type:0
  PFA_v1 g46 (.A(w11), .B(w31), .C(w37), .S(w40), .P(w30), .G(w29));   //: @(-838, 403) /sz:(126, 115) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>5 Bo0<0 Bo1<0 Bo2<0 ]
  //: switch g57 (w41) @(-666,385) /sn:0 /w:[ 0 ] /st:1
  //: joint g150 (w81) @(-2529, 990) /w:[ 2 1 -1 4 ]
  //: switch g14 (w25) @(547,120) /sn:0 /w:[ 0 ] /st:0
  //: switch g11 (w19) @(240,118) /sn:0 /w:[ 0 ] /st:0
  //: switch g5 (w32) @(698,163) /sn:0 /w:[ 3 ] /st:1
  //: switch g84 (w50) @(-1683,588) /sn:0 /w:[ 0 ] /st:1
  led g118 (.I(w60));   //: @(-1534,624) /sn:0 /w:[ 3 ] /type:0
  led g112 (.I(w55));   //: @(-1412,778) /sn:0 /w:[ 3 ] /type:0
  //: joint g21 (w35) @(156, 187) /w:[ -1 2 4 1 ]
  //: joint g61 (w27) @(-609, 571) /w:[ 2 1 -1 4 ]
  //: joint g123 (w51) @(-1077, 811) /w:[ 2 1 -1 4 ]
  led g20 (.I(w35));   //: @(150,135) /sn:0 /w:[ 3 ] /type:0
  led g32 (.I(w10));   //: @(388,286) /sn:0 /w:[ 3 ] /type:0
  led g79 (.I(w29));   //: @(-746,579) /sn:0 /w:[ 3 ] /type:0
  //: joint g115 (w59) @(-892, 678) /w:[ -1 4 3 6 ]
  //: joint g145 (w78) @(-2311, 994) /w:[ 2 1 -1 4 ]
  led g134 (.I(w76));   //: @(-2128,1027) /sn:0 /w:[ 3 ] /type:0
  led g97 (.I(w61));   //: @(-1361,655) /sn:0 /w:[ 3 ] /type:0
  //: joint g148 (w77) @(-2182, 1001) /w:[ 2 1 -1 4 ]
  //: joint g129 (w85) @(-2048, 891) /w:[ -1 2 4 1 ]
  //: switch g15 (w26) @(604,113) /sn:0 /w:[ 0 ] /st:1
  led g89 (.I(w51));   //: @(-993,828) /sn:0 /w:[ 3 ] /type:0
  //: joint g165 (w7) @(-1945, 1017) /w:[ 2 1 -1 4 ]
  //: joint g147 (w76) @(-2151, 1031) /w:[ 2 1 -1 4 ]
  //: joint g27 (w3) @(607, 322) /w:[ 2 1 -1 4 ]
  led g160 (.I(w83));   //: @(-2402,830) /sn:0 /w:[ 3 ] /type:0
  led g62 (.I(w40));   //: @(-723,550) /sn:0 /w:[ 1 ] /type:0
  led g55 (.I(w38));   //: @(-527,438) /sn:0 /w:[ 3 ] /type:0
  PFA_v1 g88 (.A(w50), .B(w63), .C(w60), .S(w64), .P(w58), .G(w57));   //: @(-1672, 620) /sz:(126, 115) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>5 Bo0<0 Bo1<0 Bo2<0 ]
  led g140 (.I(w95));   //: @(-1913,983) /sn:0 /w:[ 0 ] /type:0
  led g139 (.I(w84));   //: @(-2229,861) /sn:0 /w:[ 3 ] /type:0
  led g135 (.I(w92));   //: @(-2113,977) /sn:0 /w:[ 0 ] /type:0
  //: switch g13 (w24) @(411,106) /sn:0 /w:[ 0 ] /st:1
  PFA_v1 g53 (.A(w45), .B(w46), .C(w39), .S(w44), .P(w13), .G(w12));   //: @(-491, 412) /sz:(126, 115) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>5 Bo0<1 Bo1<0 Bo2<0 ]

endmodule
