//: version "1.8.7"

module CarryLookahead_Logic(C3, P0, w1, G0, w0, G1, P1, P2, C2, C1, G3, Cin, G2);
//: interface  /sz:(328, 96) /bd:[ Ti0>G0(286/328) Ti1>P0(267/328) Ti2>G1(210/328) Ti3>P1(189/328) Ti4>G2(139/328) Ti5>P2(117/328) Ti6>G3(55/328) Ti7>P3(28/328) Ri0>Cin(46/96) To0<C3(86/328) To1<C2(159/328) To2<C1(228/328) Lo0<Cout(39/96) ]
input G2;    //: /sn:0 /dp:1 {0}(559,261)(537,261)(537,282)(527,282)(527,313)(49,313){1}
input P1;    //: /sn:0 /dp:1 {0}(336,157)(326,157)(326,178)(316,178)(316,230)(53,230){1}
input w0;    //: /sn:0 {0}(40,343)(48,343)(48,323)(599,323)(599,302)(617,302){1}
output C3;    //: /sn:0 /dp:1 {0}(580,259)(592,259)(592,278)(595,278){1}
//: {2}(599,278)(618,278)(618,269)(622,269){3}
//: {4}(597,280)(597,297)(617,297){5}
input G0;    //: /sn:0 {0}(72,169)(254,169)(254,139)(264,139)(264,129){1}
//: {2}(266,127)(270,127){3}
//: {4}(262,127)(258,127){5}
output C2;    //: /sn:0 /dp:1 {0}(417,169)(429,169)(429,178)(432,178){1}
//: {2}(436,178)(454,178)(454,177)(456,177){3}
//: {4}(434,180)(434,246)(466,246){5}
output w1;    //: /sn:0 {0}(699,317)(734,317)(734,333)(758,333){1}
input Cin;    //: /sn:0 {0}(85,65)(97,65){1}
//: {2}(101,65)(108,65){3}
//: {4}(99,67)(99,82)(151,82){5}
input G1;    //: /sn:0 /dp:1 {0}(396,171)(381,171)(381,180)(371,180)(371,249)(51,249){1}
input G3;    //: /sn:0 {0}(30,372)(681,372)(681,339)(669,339)(669,319)(678,319){1}
output C1;    //: /sn:0 /dp:1 {0}(291,125)(295,125)(295,112)(304,112)(304,127)(314,127){1}
//: {2}(318,127)(349,127)(349,125)(352,125){3}
//: {4}(316,129)(316,152)(336,152){5}
input P0;    //: /sn:0 {0}(72,145)(132,145)(132,87)(151,87){1}
input P2;    //: /sn:0 /dp:1 {0}(466,251)(462,251)(462,277)(452,277)(452,284)(50,284){1}
wire w4;    //: /sn:0 {0}(357,155)(364,155)(364,166)(396,166){1}
wire w3;    //: /sn:0 {0}(487,249)(514,249)(514,256)(559,256){1}
wire w2;    //: /sn:0 {0}(638,300)(668,300)(668,314)(678,314){1}
wire w5;    //: /sn:0 {0}(258,124)(258,118){1}
//: {2}(260,116)(265,116)(265,122)(270,122){3}
//: {4}(258,114)(258,85)(172,85){5}
//: enddecls

  and g4 (.I0(Cin), .I1(P0), .Z(w5));   //: @(162,85) /sn:0 /tech:unit /w:[ 5 1 5 ]
  and g8 (.I0(C1), .I1(P1), .Z(w4));   //: @(347,155) /sn:0 /tech:unit /w:[ 5 0 0 ]
  or g3 (.I0(w5), .I1(G0), .Z(C1));   //: @(281,125) /sn:0 /tech:unit /w:[ 3 3 0 ]
  or g16 (.I0(w3), .I1(G2), .Z(C3));   //: @(570,259) /sn:0 /tech:unit /w:[ 1 0 0 ]
  //: output g17 (C3) @(619,269) /sn:0 /w:[ 3 ]
  //: joint g26 (C1) @(316, 127) /w:[ 2 -1 1 4 ]
  //: input g2 (P0) @(70,145) /sn:0 /w:[ 0 ]
  //: output g23 (w1) @(755,333) /sn:0 /w:[ 1 ]
  //: input g1 (G0) @(70,169) /sn:0 /w:[ 0 ]
  //: joint g24 (Cin) @(99, 65) /w:[ 2 -1 1 4 ]
  //: input g18 (w0) @(38,343) /sn:0 /w:[ 0 ]
  //: joint g25 (G0) @(264, 127) /w:[ 2 -1 4 1 ]
  or g10 (.I0(w4), .I1(G1), .Z(C2));   //: @(407,169) /sn:0 /tech:unit /w:[ 1 0 0 ]
  //: input g6 (G1) @(49,249) /sn:0 /w:[ 1 ]
  //: input g7 (P1) @(51,230) /sn:0 /w:[ 1 ]
  //: joint g9 (w5) @(258, 116) /w:[ 2 4 -1 1 ]
  or g22 (.I0(w2), .I1(G3), .Z(w1));   //: @(689,317) /sn:0 /tech:unit /w:[ 1 1 0 ]
  //: input g12 (P2) @(48,284) /sn:0 /w:[ 1 ]
  //: joint g28 (C3) @(597, 278) /w:[ 2 -1 1 4 ]
  //: output g11 (C2) @(453,177) /sn:0 /w:[ 3 ]
  //: output g5 (C1) @(349,125) /sn:0 /w:[ 3 ]
  and g14 (.I0(C2), .I1(P2), .Z(w3));   //: @(477,249) /sn:0 /tech:unit /w:[ 5 0 0 ]
  //: input g19 (G3) @(28,372) /sn:0 /w:[ 0 ]
  and g20 (.I0(C3), .I1(w0), .Z(w2));   //: @(628,300) /sn:0 /tech:unit /w:[ 5 1 0 ]
  //: input g0 (Cin) @(83,65) /sn:0 /w:[ 0 ]
  //: joint g27 (C2) @(434, 178) /w:[ 2 -1 1 4 ]
  //: input g13 (G2) @(47,313) /sn:0 /w:[ 1 ]

endmodule

module main;    //: root_module
wire w6;    //: /sn:0 {0}(306,98)(306,108){1}
wire w7;    //: /sn:0 {0}(284,98)(284,108){1}
wire w4;    //: /sn:0 {0}(377,98)(377,108){1}
wire w3;    //: /sn:0 {0}(434,98)(434,108){1}
wire w0;    //: /sn:0 {0}(506,155)(496,155){1}
wire w12;    //: /sn:0 {0}(395,98)(395,108){1}
wire w10;    //: /sn:0 {0}(253,98)(253,108){1}
wire w1;    //: /sn:0 {0}(156,148)(166,148){1}
wire w8;    //: /sn:0 {0}(222,98)(222,108){1}
wire w11;    //: /sn:0 {0}(326,98)(326,108){1}
wire w2;    //: /sn:0 {0}(453,98)(453,108){1}
wire w5;    //: /sn:0 {0}(356,98)(356,108){1}
wire w9;    //: /sn:0 {0}(195,98)(195,108){1}
//: enddecls

  CarryLookahead_Logic g0 (.P3(w9), .G3(w8), .P2(w7), .G2(w6), .P1(w5), .G1(w4), .P0(w3), .G0(w2), .Cin(w0), .C1(w12), .C2(w11), .C3(w10), .Cout(w1));   //: @(167, 109) /sz:(328, 96) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Ti3>1 Ti4>1 Ti5>1 Ti6>1 Ti7>1 Ri0>1 To0<1 To1<1 To2<1 Lo0<1 ]

endmodule
